
module MIPS ( clk, rst, pc_rom, inst_rom, ram_size, ram_read, ram_write, 
        ram_data, ram_word, ram_adr );
  output [31:0] pc_rom;
  input [31:0] inst_rom;
  output [1:0] ram_size;
  output [31:0] ram_data;
  input [31:0] ram_word;
  output [31:0] ram_adr;
  input clk, rst;
  output ram_read, ram_write;
  wire   reg_write, \wb_WB[0] , \instruction_fetch/n87 ,
         \instruction_fetch/n86 , \instruction_fetch/mux/N14 ,
         \instruction_fetch/mux/N13 , \instruction_decode/N22 ,
         \instruction_decode/N21 , \instruction_decode/N20 ,
         \instruction_decode/N19 , \instruction_decode/N18 ,
         \instruction_decode/N17 , \instruction_decode/N16 ,
         \instruction_decode/N15 , \instruction_decode/N14 ,
         \instruction_decode/N13 , \instruction_decode/N12 ,
         \instruction_decode/N11 , \instruction_decode/old_wb[1] ,
         \instruction_decode/reg_MAPP/n1276 ,
         \instruction_decode/reg_MAPP/n1275 ,
         \instruction_decode/reg_MAPP/n1274 ,
         \instruction_decode/reg_MAPP/n1273 ,
         \instruction_decode/reg_MAPP/n1272 ,
         \instruction_decode/reg_MAPP/n1271 ,
         \instruction_decode/reg_MAPP/n1270 ,
         \instruction_decode/reg_MAPP/n1269 ,
         \instruction_decode/reg_MAPP/n1268 ,
         \instruction_decode/reg_MAPP/n1267 ,
         \instruction_decode/reg_MAPP/n1266 ,
         \instruction_decode/reg_MAPP/n1265 ,
         \instruction_decode/reg_MAPP/n1264 ,
         \instruction_decode/reg_MAPP/n1263 ,
         \instruction_decode/reg_MAPP/n1262 ,
         \instruction_decode/reg_MAPP/n1261 ,
         \instruction_decode/reg_MAPP/n1260 ,
         \instruction_decode/reg_MAPP/n1259 ,
         \instruction_decode/reg_MAPP/n1258 ,
         \instruction_decode/reg_MAPP/n1257 ,
         \instruction_decode/reg_MAPP/n1256 ,
         \instruction_decode/reg_MAPP/n1255 ,
         \instruction_decode/reg_MAPP/n1254 ,
         \instruction_decode/reg_MAPP/n1253 ,
         \instruction_decode/reg_MAPP/n1252 ,
         \instruction_decode/reg_MAPP/n1251 ,
         \instruction_decode/reg_MAPP/n1250 ,
         \instruction_decode/reg_MAPP/n1249 ,
         \instruction_decode/reg_MAPP/n1248 ,
         \instruction_decode/reg_MAPP/n1247 ,
         \instruction_decode/reg_MAPP/n1246 ,
         \instruction_decode/reg_MAPP/n1245 ,
         \instruction_decode/reg_MAPP/n3641 ,
         \instruction_decode/hazard_unit/n5 , \execute/n459 , \execute/n453 ,
         \execute/n434 , \execute/n433 , \execute/n432 , \execute/n431 ,
         \execute/n430 , \execute/alu/sll_175/ML_int[5][16] ,
         \execute/alu/sll_175/ML_int[5][17] ,
         \execute/alu/sll_175/ML_int[5][19] ,
         \execute/alu/sll_175/ML_int[5][20] ,
         \execute/alu/sll_175/ML_int[5][21] ,
         \execute/alu/sll_175/ML_int[5][23] ,
         \execute/alu/sll_175/ML_int[5][24] ,
         \execute/alu/sll_175/ML_int[5][25] ,
         \execute/alu/sll_175/ML_int[5][26] ,
         \execute/alu/sll_175/ML_int[5][27] ,
         \execute/alu/sll_175/ML_int[5][28] ,
         \execute/alu/sll_175/ML_int[5][29] ,
         \execute/alu/sll_175/ML_int[5][30] ,
         \execute/alu/sll_175/ML_int[4][8] ,
         \execute/alu/sll_175/ML_int[4][9] ,
         \execute/alu/sll_175/ML_int[4][10] ,
         \execute/alu/sll_175/ML_int[4][11] ,
         \execute/alu/sll_175/ML_int[4][12] ,
         \execute/alu/sll_175/ML_int[4][13] ,
         \execute/alu/sll_175/ML_int[4][14] ,
         \execute/alu/sll_175/ML_int[4][17] ,
         \execute/alu/sll_175/ML_int[4][21] ,
         \execute/alu/sll_175/ML_int[4][23] ,
         \execute/alu/sll_175/ML_int[4][24] ,
         \execute/alu/sll_175/ML_int[4][25] ,
         \execute/alu/sll_175/ML_int[4][26] ,
         \execute/alu/sll_175/ML_int[4][27] ,
         \execute/alu/sll_175/ML_int[4][28] ,
         \execute/alu/sll_175/ML_int[4][29] ,
         \execute/alu/sll_175/ML_int[4][30] ,
         \execute/alu/sll_175/ML_int[3][4] ,
         \execute/alu/sll_175/ML_int[3][5] ,
         \execute/alu/sll_175/ML_int[3][6] ,
         \execute/alu/sll_175/ML_int[3][7] ,
         \execute/alu/sll_175/ML_int[3][8] ,
         \execute/alu/sll_175/ML_int[3][9] ,
         \execute/alu/sll_175/ML_int[3][10] ,
         \execute/alu/sll_175/ML_int[3][11] ,
         \execute/alu/sll_175/ML_int[3][12] ,
         \execute/alu/sll_175/ML_int[3][13] ,
         \execute/alu/sll_175/ML_int[3][14] ,
         \execute/alu/sll_175/ML_int[3][15] ,
         \execute/alu/sll_175/ML_int[3][16] ,
         \execute/alu/sll_175/ML_int[3][17] ,
         \execute/alu/sll_175/ML_int[3][18] ,
         \execute/alu/sll_175/ML_int[3][19] ,
         \execute/alu/sll_175/ML_int[3][20] ,
         \execute/alu/sll_175/ML_int[3][21] ,
         \execute/alu/sll_175/ML_int[3][22] ,
         \execute/alu/sll_175/ML_int[3][23] ,
         \execute/alu/sll_175/ML_int[3][24] ,
         \execute/alu/sll_175/ML_int[3][25] ,
         \execute/alu/sll_175/ML_int[3][26] ,
         \execute/alu/sll_175/ML_int[3][27] ,
         \execute/alu/sll_175/ML_int[3][28] ,
         \execute/alu/sll_175/ML_int[3][29] ,
         \execute/alu/sll_175/ML_int[3][30] ,
         \execute/alu/sll_175/ML_int[2][0] ,
         \execute/alu/sll_175/ML_int[2][2] ,
         \execute/alu/sll_175/ML_int[2][3] ,
         \execute/alu/sll_175/ML_int[2][4] ,
         \execute/alu/sll_175/ML_int[2][5] ,
         \execute/alu/sll_175/ML_int[2][6] ,
         \execute/alu/sll_175/ML_int[2][7] ,
         \execute/alu/sll_175/ML_int[2][8] ,
         \execute/alu/sll_175/ML_int[2][9] ,
         \execute/alu/sll_175/ML_int[2][10] ,
         \execute/alu/sll_175/ML_int[2][11] ,
         \execute/alu/sll_175/ML_int[2][12] ,
         \execute/alu/sll_175/ML_int[2][13] ,
         \execute/alu/sll_175/ML_int[2][14] ,
         \execute/alu/sll_175/ML_int[2][15] ,
         \execute/alu/sll_175/ML_int[2][16] ,
         \execute/alu/sll_175/ML_int[2][17] ,
         \execute/alu/sll_175/ML_int[2][18] ,
         \execute/alu/sll_175/ML_int[2][19] ,
         \execute/alu/sll_175/ML_int[2][20] ,
         \execute/alu/sll_175/ML_int[2][21] ,
         \execute/alu/sll_175/ML_int[2][22] ,
         \execute/alu/sll_175/ML_int[2][23] ,
         \execute/alu/sll_175/ML_int[2][24] ,
         \execute/alu/sll_175/ML_int[2][25] ,
         \execute/alu/sll_175/ML_int[2][26] ,
         \execute/alu/sll_175/ML_int[2][27] ,
         \execute/alu/sll_175/ML_int[2][28] ,
         \execute/alu/sll_175/ML_int[2][29] ,
         \execute/alu/sll_175/ML_int[2][30] ,
         \execute/alu/sll_175/ML_int[2][31] ,
         \execute/alu/sll_175/ML_int[1][1] ,
         \execute/alu/sll_175/ML_int[1][2] ,
         \execute/alu/sll_175/ML_int[1][3] ,
         \execute/alu/sll_175/ML_int[1][4] ,
         \execute/alu/sll_175/ML_int[1][5] ,
         \execute/alu/sll_175/ML_int[1][6] ,
         \execute/alu/sll_175/ML_int[1][7] ,
         \execute/alu/sll_175/ML_int[1][8] ,
         \execute/alu/sll_175/ML_int[1][9] ,
         \execute/alu/sll_175/ML_int[1][10] ,
         \execute/alu/sll_175/ML_int[1][11] ,
         \execute/alu/sll_175/ML_int[1][12] ,
         \execute/alu/sll_175/ML_int[1][13] ,
         \execute/alu/sll_175/ML_int[1][14] ,
         \execute/alu/sll_175/ML_int[1][15] ,
         \execute/alu/sll_175/ML_int[1][16] ,
         \execute/alu/sll_175/ML_int[1][17] ,
         \execute/alu/sll_175/ML_int[1][18] ,
         \execute/alu/sll_175/ML_int[1][19] ,
         \execute/alu/sll_175/ML_int[1][20] ,
         \execute/alu/sll_175/ML_int[1][21] ,
         \execute/alu/sll_175/ML_int[1][22] ,
         \execute/alu/sll_175/ML_int[1][23] ,
         \execute/alu/sll_175/ML_int[1][24] ,
         \execute/alu/sll_175/ML_int[1][25] ,
         \execute/alu/sll_175/ML_int[1][26] ,
         \execute/alu/sll_175/ML_int[1][27] ,
         \execute/alu/sll_175/ML_int[1][28] ,
         \execute/alu/sll_175/ML_int[1][29] ,
         \execute/alu/sll_175/ML_int[1][30] ,
         \execute/alu/sll_175/ML_int[1][31] ,
         \execute/alu/sll_175/temp_int_SH[0] ,
         \execute/alu/sll_175/temp_int_SH[1] ,
         \execute/alu/sll_175/temp_int_SH[2] ,
         \execute/alu/sll_175/temp_int_SH[3] ,
         \execute/alu/sll_175/temp_int_SH[4] , n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1185, n1187, n1211, n1214, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1257, n1258, n1259, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1338, n1339, n1340, n1341, n1342, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1433, n1434, n1435, n1436, n1437, n1439, n1440, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1465,
         n1467, n1468, n1470, n1471, n1472, n1473, n1476, n1478, n1481, n1484,
         n1485, n1486, n1489, n1490, n1491, n1492, n1493, n1494, n1728, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1952, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2036, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4575, n4576, n4577, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4714, n4718, n4722, n4726, n4730, n4734, n4738, n4742, n4746,
         n4750, n4754, n4758, n4762, n4766, n4770, n4774, n4778, n4782, n4786,
         n4790, n4794, n4798, n4802, n4806, n4810, n4814, n4818, n4822, n4826,
         n4830, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5308, n5309, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5356, n5358, n5359, n5360, n5362,
         n5363, n5364, n5368, n5370, n5371, n5372, n5376, n5378, n5379, n5380,
         n5384, n5386, n5387, n5388, n5392, n5394, n5395, n5396, n5400, n5402,
         n5403, n5404, n5408, n5410, n5411, n5412, n5416, n5418, n5419, n5420,
         n5424, n5426, n5427, n5428, n5432, n5434, n5435, n5436, n5440, n5442,
         n5443, n5444, n5446, n5447, n5448, n5452, n5454, n5455, n5456, n5460,
         n5462, n5463, n5464, n5468, n5470, n5471, n5472, n5476, n5478, n5479,
         n5480, n5484, n5486, n5487, n5488, n5492, n5494, n5495, n5496, n5500,
         n5502, n5503, n5504, n5508, n5510, n5511, n5512, n5516, n5518, n5519,
         n5520, n5524, n5526, n5527, n5528, n5532, n5534, n5535, n5536, n5540,
         n5542, n5543, n5544, n5548, n5550, n5551, n5552, n5556, n5558, n5559,
         n5560, n5564, n5566, n5567, n5568, n5572, n5574, n5575, n5576, n5580,
         n5582, n5583, n5584, n5588, n5590, n5591, n5592, n5596, n5598, n5599,
         n5600, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5617, n5619, n5620, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5694, n5695, n5696, n5697, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994;
  wire   [31:0] pc_branch;
  wire   [31:0] pc_out;
  wire   [31:0] inst_out;
  wire   [4:0] write_register;
  wire   [31:0] write_data_reg;
  wire   [4:0] rs;
  wire   [4:0] rt;
  wire   [31:0] data_1;
  wire   [31:0] data_2;
  wire   [31:0] pc_ex;
  wire   [4:0] write_register_ex;
  wire   [1:0] wb_MEM;
  wire   [31:0] \instruction_fetch/pc_4 ;
  wire   [4:0] \instruction_decode/old_rd ;
  wire   [5:0] \instruction_decode/old_ex ;
  wire   [3:0] \instruction_decode/old_m ;
  wire   [31:0] \instruction_decode/old_data_2 ;
  wire   [31:0] \instruction_decode/old_data_1 ;
  wire   [15:1] \instruction_decode/add_358/carry ;
  wire   [31:0] \execute/op_21 ;
  wire   [31:0] \execute/old_res ;
  assign pc_rom[2] = \instruction_fetch/n87 ;
  assign pc_rom[3] = \instruction_fetch/n86 ;
  assign pc_rom[1] = \instruction_fetch/mux/N14 ;
  assign pc_rom[0] = \instruction_fetch/mux/N13 ;

  DF3 \instruction_fetch/pc_out_reg[0]  ( .D(\instruction_fetch/mux/N13 ), .C(
        clk), .Q(pc_out[0]), .QN(n5709) );
  DF3 \instruction_fetch/pc_out_reg[1]  ( .D(\instruction_fetch/mux/N14 ), .C(
        clk), .Q(pc_out[1]), .QN(n5708) );
  DF3 \instruction_fetch/pc_out_reg[2]  ( .D(\instruction_fetch/n87 ), .C(clk), 
        .Q(pc_out[2]), .QN(n6080) );
  DF3 \instruction_fetch/pc_out_reg[3]  ( .D(\instruction_fetch/n86 ), .C(clk), 
        .Q(pc_out[3]) );
  DF3 \instruction_fetch/pc_out_reg[4]  ( .D(pc_rom[4]), .C(clk), .Q(pc_out[4]) );
  DF3 \instruction_fetch/pc_out_reg[5]  ( .D(pc_rom[5]), .C(clk), .Q(pc_out[5]) );
  DF3 \instruction_fetch/pc_out_reg[6]  ( .D(pc_rom[6]), .C(clk), .Q(pc_out[6]) );
  DF3 \instruction_fetch/pc_out_reg[7]  ( .D(pc_rom[7]), .C(clk), .Q(pc_out[7]) );
  DF3 \instruction_fetch/pc_out_reg[8]  ( .D(pc_rom[8]), .C(clk), .Q(pc_out[8]) );
  DF3 \instruction_fetch/pc_out_reg[9]  ( .D(pc_rom[9]), .C(clk), .Q(pc_out[9]) );
  DF3 \instruction_fetch/pc_out_reg[10]  ( .D(pc_rom[10]), .C(clk), .Q(
        pc_out[10]) );
  DF3 \instruction_fetch/pc_out_reg[11]  ( .D(pc_rom[11]), .C(clk), .Q(
        pc_out[11]) );
  DF3 \instruction_fetch/pc_out_reg[12]  ( .D(pc_rom[12]), .C(clk), .Q(
        pc_out[12]) );
  DF3 \instruction_fetch/pc_out_reg[13]  ( .D(pc_rom[13]), .C(clk), .Q(
        pc_out[13]) );
  DF3 \instruction_fetch/pc_out_reg[14]  ( .D(pc_rom[14]), .C(clk), .Q(
        pc_out[14]) );
  DF3 \instruction_fetch/pc_out_reg[15]  ( .D(pc_rom[15]), .C(clk), .Q(
        pc_out[15]), .QN(n6263) );
  DF3 \instruction_fetch/pc_out_reg[16]  ( .D(pc_rom[16]), .C(clk), .Q(
        pc_out[16]) );
  DF3 \instruction_fetch/pc_out_reg[17]  ( .D(pc_rom[17]), .C(clk), .Q(
        pc_out[17]), .QN(n5707) );
  DF3 \instruction_fetch/pc_out_reg[18]  ( .D(pc_rom[18]), .C(clk), .Q(
        pc_out[18]) );
  DF3 \instruction_fetch/pc_out_reg[19]  ( .D(pc_rom[19]), .C(clk), .Q(
        pc_out[19]), .QN(n5706) );
  DF3 \instruction_fetch/pc_out_reg[20]  ( .D(pc_rom[20]), .C(clk), .Q(
        pc_out[20]) );
  DF3 \instruction_fetch/pc_out_reg[21]  ( .D(pc_rom[21]), .C(clk), .Q(
        pc_out[21]), .QN(n5705) );
  DF3 \instruction_fetch/pc_out_reg[22]  ( .D(pc_rom[22]), .C(clk), .Q(
        pc_out[22]) );
  DF3 \instruction_fetch/pc_out_reg[23]  ( .D(pc_rom[23]), .C(clk), .Q(
        pc_out[23]), .QN(n5704) );
  DF3 \instruction_fetch/pc_out_reg[24]  ( .D(pc_rom[24]), .C(clk), .Q(
        pc_out[24]) );
  DF3 \instruction_fetch/pc_out_reg[25]  ( .D(pc_rom[25]), .C(clk), .Q(
        pc_out[25]), .QN(n5703) );
  DF3 \instruction_fetch/pc_out_reg[26]  ( .D(pc_rom[26]), .C(clk), .Q(
        pc_out[26]) );
  DF3 \instruction_fetch/pc_out_reg[27]  ( .D(pc_rom[27]), .C(clk), .Q(
        pc_out[27]), .QN(n5702) );
  DF3 \instruction_fetch/pc_out_reg[28]  ( .D(pc_rom[28]), .C(clk), .Q(
        pc_branch[28]), .QN(n6272) );
  DF3 \instruction_fetch/pc_out_reg[29]  ( .D(pc_rom[29]), .C(clk), .Q(
        pc_branch[29]), .QN(n4575) );
  DF3 \instruction_fetch/pc_out_reg[30]  ( .D(pc_rom[30]), .C(clk), .Q(
        pc_branch[30]), .QN(n4579) );
  DF3 \instruction_fetch/pc_out_reg[31]  ( .D(pc_rom[31]), .C(clk), .Q(
        pc_branch[31]), .QN(n6276) );
  DF3 \instruction_decode/pc_ex_reg[0]  ( .D(pc_out[0]), .C(clk), .Q(pc_ex[0])
         );
  DF3 \instruction_decode/pc_ex_reg[1]  ( .D(pc_out[1]), .C(clk), .Q(pc_ex[1])
         );
  DF3 \instruction_decode/pc_ex_reg[2]  ( .D(pc_out[2]), .C(clk), .Q(pc_ex[2])
         );
  DF3 \instruction_decode/pc_ex_reg[3]  ( .D(pc_out[3]), .C(clk), .Q(pc_ex[3])
         );
  DF3 \instruction_decode/pc_ex_reg[4]  ( .D(pc_out[4]), .C(clk), .Q(pc_ex[4])
         );
  DF3 \instruction_decode/pc_ex_reg[5]  ( .D(pc_out[5]), .C(clk), .Q(pc_ex[5])
         );
  DF3 \instruction_decode/pc_ex_reg[6]  ( .D(pc_out[6]), .C(clk), .Q(pc_ex[6])
         );
  DF3 \instruction_decode/pc_ex_reg[7]  ( .D(pc_out[7]), .C(clk), .Q(pc_ex[7])
         );
  DF3 \instruction_decode/pc_ex_reg[8]  ( .D(pc_out[8]), .C(clk), .Q(pc_ex[8])
         );
  DF3 \instruction_decode/pc_ex_reg[9]  ( .D(pc_out[9]), .C(clk), .Q(pc_ex[9])
         );
  DF3 \instruction_decode/pc_ex_reg[10]  ( .D(pc_out[10]), .C(clk), .Q(
        pc_ex[10]) );
  DF3 \instruction_decode/pc_ex_reg[11]  ( .D(pc_out[11]), .C(clk), .Q(
        pc_ex[11]) );
  DF3 \instruction_decode/pc_ex_reg[12]  ( .D(pc_out[12]), .C(clk), .Q(
        pc_ex[12]) );
  DF3 \instruction_decode/pc_ex_reg[13]  ( .D(pc_out[13]), .C(clk), .Q(
        pc_ex[13]) );
  DF3 \instruction_decode/pc_ex_reg[14]  ( .D(pc_out[14]), .C(clk), .Q(
        pc_ex[14]) );
  DF3 \instruction_decode/pc_ex_reg[15]  ( .D(pc_out[15]), .C(clk), .Q(
        pc_ex[15]) );
  DF3 \instruction_decode/pc_ex_reg[16]  ( .D(pc_out[16]), .C(clk), .Q(
        pc_ex[16]) );
  DF3 \instruction_decode/pc_ex_reg[17]  ( .D(pc_out[17]), .C(clk), .Q(
        pc_ex[17]) );
  DF3 \instruction_decode/pc_ex_reg[18]  ( .D(pc_out[18]), .C(clk), .Q(
        pc_ex[18]) );
  DF3 \instruction_decode/pc_ex_reg[19]  ( .D(pc_out[19]), .C(clk), .Q(
        pc_ex[19]) );
  DF3 \instruction_decode/pc_ex_reg[20]  ( .D(pc_out[20]), .C(clk), .Q(
        pc_ex[20]) );
  DF3 \instruction_decode/pc_ex_reg[21]  ( .D(pc_out[21]), .C(clk), .Q(
        pc_ex[21]) );
  DF3 \instruction_decode/pc_ex_reg[22]  ( .D(pc_out[22]), .C(clk), .Q(
        pc_ex[22]) );
  DF3 \instruction_decode/pc_ex_reg[23]  ( .D(pc_out[23]), .C(clk), .Q(
        pc_ex[23]) );
  DF3 \instruction_decode/pc_ex_reg[24]  ( .D(pc_out[24]), .C(clk), .Q(
        pc_ex[24]) );
  DF3 \instruction_decode/pc_ex_reg[25]  ( .D(pc_out[25]), .C(clk), .Q(
        pc_ex[25]) );
  DF3 \instruction_decode/pc_ex_reg[26]  ( .D(pc_out[26]), .C(clk), .Q(
        pc_ex[26]) );
  DF3 \instruction_decode/pc_ex_reg[27]  ( .D(pc_out[27]), .C(clk), .Q(
        pc_ex[27]) );
  DF3 \instruction_decode/pc_ex_reg[28]  ( .D(pc_branch[28]), .C(clk), .Q(
        pc_ex[28]) );
  DF3 \instruction_decode/pc_ex_reg[29]  ( .D(pc_branch[29]), .C(clk), .Q(
        pc_ex[29]) );
  DF3 \instruction_decode/pc_ex_reg[30]  ( .D(pc_branch[30]), .C(clk), .Q(
        pc_ex[30]), .QN(n5612) );
  DF3 \instruction_decode/pc_ex_reg[31]  ( .D(pc_branch[31]), .C(clk), .Q(
        pc_ex[31]) );
  DF3 \instruction_decode/data_2_reg[0]  ( .D(
        \instruction_decode/old_data_2 [0]), .C(clk), .Q(data_2[0]) );
  DF3 \instruction_decode/data_2_reg[1]  ( .D(
        \instruction_decode/old_data_2 [1]), .C(clk), .Q(data_2[1]) );
  DF3 \instruction_decode/data_2_reg[2]  ( .D(
        \instruction_decode/old_data_2 [2]), .C(clk), .Q(data_2[2]) );
  DF3 \instruction_decode/data_2_reg[3]  ( .D(
        \instruction_decode/old_data_2 [3]), .C(clk), .Q(data_2[3]) );
  DF3 \instruction_decode/data_2_reg[4]  ( .D(
        \instruction_decode/old_data_2 [4]), .C(clk), .Q(data_2[4]) );
  DF3 \instruction_decode/data_2_reg[5]  ( .D(
        \instruction_decode/old_data_2 [5]), .C(clk), .Q(data_2[5]) );
  DF3 \instruction_decode/data_2_reg[6]  ( .D(
        \instruction_decode/old_data_2 [6]), .C(clk), .Q(data_2[6]) );
  DF3 \instruction_decode/data_2_reg[7]  ( .D(
        \instruction_decode/old_data_2 [7]), .C(clk), .Q(data_2[7]) );
  DF3 \instruction_decode/data_2_reg[8]  ( .D(
        \instruction_decode/old_data_2 [8]), .C(clk), .Q(data_2[8]) );
  DF3 \instruction_decode/data_2_reg[9]  ( .D(
        \instruction_decode/old_data_2 [9]), .C(clk), .Q(data_2[9]) );
  DF3 \instruction_decode/data_2_reg[10]  ( .D(
        \instruction_decode/old_data_2 [10]), .C(clk), .Q(data_2[10]) );
  DF3 \instruction_decode/data_2_reg[11]  ( .D(
        \instruction_decode/old_data_2 [11]), .C(clk), .Q(data_2[11]) );
  DF3 \instruction_decode/data_2_reg[12]  ( .D(
        \instruction_decode/old_data_2 [12]), .C(clk), .Q(data_2[12]) );
  DF3 \instruction_decode/data_2_reg[13]  ( .D(
        \instruction_decode/old_data_2 [13]), .C(clk), .Q(data_2[13]) );
  DF3 \instruction_decode/data_2_reg[14]  ( .D(
        \instruction_decode/old_data_2 [14]), .C(clk), .Q(data_2[14]) );
  DF3 \instruction_decode/data_2_reg[15]  ( .D(
        \instruction_decode/old_data_2 [15]), .C(clk), .Q(data_2[15]) );
  DF3 \instruction_decode/data_2_reg[16]  ( .D(
        \instruction_decode/old_data_2 [16]), .C(clk), .Q(data_2[16]) );
  DF3 \instruction_decode/data_2_reg[17]  ( .D(
        \instruction_decode/old_data_2 [17]), .C(clk), .Q(data_2[17]) );
  DF3 \instruction_decode/data_2_reg[18]  ( .D(
        \instruction_decode/old_data_2 [18]), .C(clk), .Q(data_2[18]) );
  DF3 \instruction_decode/data_2_reg[19]  ( .D(
        \instruction_decode/old_data_2 [19]), .C(clk), .Q(data_2[19]) );
  DF3 \instruction_decode/data_2_reg[20]  ( .D(
        \instruction_decode/old_data_2 [20]), .C(clk), .Q(data_2[20]) );
  DF3 \instruction_decode/data_2_reg[21]  ( .D(
        \instruction_decode/old_data_2 [21]), .C(clk), .Q(data_2[21]) );
  DF3 \instruction_decode/data_2_reg[22]  ( .D(
        \instruction_decode/old_data_2 [22]), .C(clk), .Q(data_2[22]) );
  DF3 \instruction_decode/data_2_reg[23]  ( .D(
        \instruction_decode/old_data_2 [23]), .C(clk), .Q(data_2[23]) );
  DF3 \instruction_decode/data_2_reg[24]  ( .D(
        \instruction_decode/old_data_2 [24]), .C(clk), .Q(data_2[24]) );
  DF3 \instruction_decode/data_2_reg[25]  ( .D(
        \instruction_decode/old_data_2 [25]), .C(clk), .Q(data_2[25]) );
  DF3 \instruction_decode/data_2_reg[26]  ( .D(
        \instruction_decode/old_data_2 [26]), .C(clk), .Q(data_2[26]) );
  DF3 \instruction_decode/data_2_reg[27]  ( .D(
        \instruction_decode/old_data_2 [27]), .C(clk), .Q(data_2[27]) );
  DF3 \instruction_decode/data_2_reg[28]  ( .D(
        \instruction_decode/old_data_2 [28]), .C(clk), .Q(data_2[28]) );
  DF3 \instruction_decode/data_2_reg[29]  ( .D(
        \instruction_decode/old_data_2 [29]), .C(clk), .Q(data_2[29]) );
  DF3 \instruction_decode/data_2_reg[30]  ( .D(
        \instruction_decode/old_data_2 [30]), .C(clk), .Q(data_2[30]) );
  DF3 \instruction_decode/data_2_reg[31]  ( .D(
        \instruction_decode/old_data_2 [31]), .C(clk), .Q(data_2[31]) );
  DF3 \instruction_decode/data_1_reg[0]  ( .D(
        \instruction_decode/old_data_1 [0]), .C(clk), .Q(data_1[0]) );
  DF3 \instruction_decode/data_1_reg[1]  ( .D(
        \instruction_decode/old_data_1 [1]), .C(clk), .Q(data_1[1]) );
  DF3 \instruction_decode/data_1_reg[2]  ( .D(
        \instruction_decode/old_data_1 [2]), .C(clk), .Q(data_1[2]) );
  DF3 \instruction_decode/data_1_reg[3]  ( .D(
        \instruction_decode/old_data_1 [3]), .C(clk), .Q(data_1[3]) );
  DF3 \instruction_decode/data_1_reg[4]  ( .D(
        \instruction_decode/old_data_1 [4]), .C(clk), .Q(data_1[4]) );
  DF3 \instruction_decode/data_1_reg[5]  ( .D(
        \instruction_decode/old_data_1 [5]), .C(clk), .Q(data_1[5]) );
  DF3 \instruction_decode/data_1_reg[6]  ( .D(
        \instruction_decode/old_data_1 [6]), .C(clk), .Q(data_1[6]) );
  DF3 \instruction_decode/data_1_reg[7]  ( .D(
        \instruction_decode/old_data_1 [7]), .C(clk), .Q(data_1[7]) );
  DF3 \instruction_decode/data_1_reg[8]  ( .D(
        \instruction_decode/old_data_1 [8]), .C(clk), .Q(data_1[8]) );
  DF3 \instruction_decode/data_1_reg[9]  ( .D(
        \instruction_decode/old_data_1 [9]), .C(clk), .Q(data_1[9]) );
  DF3 \instruction_decode/data_1_reg[10]  ( .D(
        \instruction_decode/old_data_1 [10]), .C(clk), .Q(data_1[10]) );
  DF3 \instruction_decode/data_1_reg[11]  ( .D(
        \instruction_decode/old_data_1 [11]), .C(clk), .Q(data_1[11]) );
  DF3 \instruction_decode/data_1_reg[12]  ( .D(
        \instruction_decode/old_data_1 [12]), .C(clk), .Q(data_1[12]) );
  DF3 \instruction_decode/data_1_reg[13]  ( .D(
        \instruction_decode/reg_MAPP/n3641 ), .C(clk), .Q(data_1[13]) );
  DF3 \instruction_decode/data_1_reg[14]  ( .D(
        \instruction_decode/old_data_1 [14]), .C(clk), .Q(data_1[14]) );
  DF3 \instruction_decode/data_1_reg[15]  ( .D(
        \instruction_decode/old_data_1 [15]), .C(clk), .Q(data_1[15]) );
  DF3 \instruction_decode/data_1_reg[16]  ( .D(
        \instruction_decode/old_data_1 [16]), .C(clk), .Q(data_1[16]) );
  DF3 \instruction_decode/data_1_reg[17]  ( .D(
        \instruction_decode/old_data_1 [17]), .C(clk), .Q(data_1[17]) );
  DF3 \instruction_decode/data_1_reg[18]  ( .D(
        \instruction_decode/old_data_1 [18]), .C(clk), .Q(data_1[18]) );
  DF3 \instruction_decode/data_1_reg[19]  ( .D(
        \instruction_decode/old_data_1 [19]), .C(clk), .Q(data_1[19]) );
  DF3 \instruction_decode/data_1_reg[20]  ( .D(
        \instruction_decode/old_data_1 [20]), .C(clk), .Q(data_1[20]) );
  DF3 \instruction_decode/data_1_reg[21]  ( .D(
        \instruction_decode/old_data_1 [21]), .C(clk), .Q(data_1[21]) );
  DF3 \instruction_decode/data_1_reg[22]  ( .D(
        \instruction_decode/old_data_1 [22]), .C(clk), .Q(data_1[22]) );
  DF3 \instruction_decode/data_1_reg[23]  ( .D(
        \instruction_decode/old_data_1 [23]), .C(clk), .Q(data_1[23]) );
  DF3 \instruction_decode/data_1_reg[24]  ( .D(
        \instruction_decode/old_data_1 [24]), .C(clk), .Q(data_1[24]) );
  DF3 \instruction_decode/data_1_reg[25]  ( .D(
        \instruction_decode/old_data_1 [25]), .C(clk), .Q(data_1[25]) );
  DF3 \instruction_decode/data_1_reg[26]  ( .D(
        \instruction_decode/old_data_1 [26]), .C(clk), .Q(data_1[26]) );
  DF3 \instruction_decode/data_1_reg[27]  ( .D(
        \instruction_decode/old_data_1 [27]), .C(clk), .Q(data_1[27]) );
  DF3 \instruction_decode/data_1_reg[28]  ( .D(
        \instruction_decode/old_data_1 [28]), .C(clk), .Q(data_1[28]) );
  DF3 \instruction_decode/data_1_reg[29]  ( .D(
        \instruction_decode/old_data_1 [29]), .C(clk), .Q(data_1[29]) );
  DF3 \instruction_decode/data_1_reg[30]  ( .D(
        \instruction_decode/old_data_1 [30]), .C(clk), .Q(data_1[30]) );
  DF3 \instruction_decode/data_1_reg[31]  ( .D(
        \instruction_decode/old_data_1 [31]), .C(clk), .Q(data_1[31]) );
  DF3 \instruction_decode/rd_reg[0]  ( .D(\instruction_decode/old_rd [0]), .C(
        clk), .QN(n5626) );
  DF3 \instruction_decode/rd_reg[1]  ( .D(\instruction_decode/old_rd [1]), .C(
        clk), .QN(n5625) );
  DF3 \instruction_decode/rd_reg[2]  ( .D(\instruction_decode/old_rd [2]), .C(
        clk), .QN(n5624) );
  DF3 \instruction_decode/rd_reg[3]  ( .D(\instruction_decode/old_rd [3]), .C(
        clk), .QN(n5623) );
  DF3 \instruction_decode/rd_reg[4]  ( .D(\instruction_decode/old_rd [4]), .C(
        clk), .QN(n5622) );
  DF3 \instruction_decode/wb_reg[1]  ( .D(\instruction_decode/old_wb[1] ), .C(
        clk), .QN(n5611) );
  DF3 \instruction_decode/wb_reg[0]  ( .D(n5773), .C(clk), .QN(n5608) );
  DF3 \instruction_decode/m_reg[3]  ( .D(\instruction_decode/old_m [3]), .C(
        clk), .QN(n5604) );
  DF3 \instruction_decode/m_reg[2]  ( .D(n1150), .C(clk), .QN(n5605) );
  DF3 \instruction_decode/m_reg[1]  ( .D(n5773), .C(clk), .Q(n6084), .QN(n5606) );
  DF3 \instruction_decode/m_reg[0]  ( .D(\instruction_decode/old_m [0]), .C(
        clk), .QN(n5607) );
  DF3 \instruction_decode/ex_reg[5]  ( .D(\instruction_decode/old_ex [5]), .C(
        clk), .QN(n5700) );
  DF3 \instruction_decode/ex_reg[3]  ( .D(\instruction_decode/old_ex [3]), .C(
        clk), .Q(n5999), .QN(n5699) );
  DF3 \instruction_decode/ex_reg[2]  ( .D(\instruction_decode/old_ex [2]), .C(
        clk), .Q(n6217), .QN(n5732) );
  DF3 \instruction_decode/ex_reg[1]  ( .D(\instruction_decode/old_ex [1]), .C(
        clk), .Q(n6233), .QN(n5733) );
  DF3 \instruction_decode/ex_reg[0]  ( .D(n1141), .C(clk), .Q(n5942), .QN(
        n5734) );
  DF3 \instruction_decode/rt_reg[0]  ( .D(inst_out[16]), .C(clk), .Q(rt[0]) );
  DF3 \instruction_decode/rt_reg[1]  ( .D(inst_out[17]), .C(clk), .QN(n6067)
         );
  DF3 \instruction_decode/rt_reg[2]  ( .D(inst_out[18]), .C(clk), .Q(rt[2]), 
        .QN(n6091) );
  DF3 \instruction_decode/rt_reg[3]  ( .D(inst_out[19]), .C(clk), .Q(rt[3]) );
  DF3 \instruction_decode/rt_reg[4]  ( .D(inst_out[20]), .C(clk), .Q(rt[4]), 
        .QN(n6220) );
  DF3 \instruction_decode/rs_reg[0]  ( .D(inst_out[21]), .C(clk), .Q(rs[0]) );
  DF3 \instruction_decode/rs_reg[1]  ( .D(inst_out[22]), .C(clk), .Q(rs[1]) );
  DF3 \instruction_decode/rs_reg[2]  ( .D(inst_out[23]), .C(clk), .Q(rs[2]) );
  DF3 \instruction_decode/rs_reg[3]  ( .D(inst_out[24]), .C(clk), .Q(rs[3]) );
  DF3 \instruction_decode/rs_reg[4]  ( .D(inst_out[25]), .C(clk), .Q(rs[4]) );
  DF3 \instruction_decode/imm_reg[1]  ( .D(inst_out[1]), .C(clk), .Q(n6247), 
        .QN(n5627) );
  DF3 \instruction_decode/imm_reg[2]  ( .D(inst_out[2]), .C(clk), .Q(n6232), 
        .QN(n5697) );
  DF3 \instruction_decode/imm_reg[3]  ( .D(inst_out[3]), .C(clk), .QN(n5696)
         );
  DF3 \instruction_decode/imm_reg[4]  ( .D(inst_out[4]), .C(clk), .QN(n5695)
         );
  DF3 \instruction_decode/imm_reg[5]  ( .D(inst_out[5]), .C(clk), .Q(n6246), 
        .QN(n5694) );
  DF3 \instruction_decode/imm_reg[6]  ( .D(inst_out[6]), .C(clk), .Q(n5944) );
  DF3 \instruction_decode/imm_reg[8]  ( .D(inst_out[8]), .C(clk), .Q(n6074) );
  DF3 \instruction_decode/imm_reg[9]  ( .D(inst_out[9]), .C(clk), .Q(n6075) );
  DF3 \instruction_decode/imm_reg[10]  ( .D(inst_out[10]), .C(clk), .Q(n6073)
         );
  DF3 \instruction_decode/imm_reg[11]  ( .D(inst_out[11]), .C(clk), .QN(n5617)
         );
  DF3 \instruction_decode/imm_reg[12]  ( .D(inst_out[12]), .C(clk), .QN(n5620)
         );
  DF3 \instruction_decode/imm_reg[13]  ( .D(inst_out[13]), .C(clk), .QN(n5610)
         );
  DF3 \instruction_decode/imm_reg[14]  ( .D(inst_out[14]), .C(clk), .QN(n5609)
         );
  DF3 \instruction_decode/imm_reg[15]  ( .D(inst_out[15]), .C(clk), .QN(n5619)
         );
  ADD32 \instruction_decode/add_358/U1_3  ( .A(pc_out[3]), .B(inst_out[1]), 
        .CI(\instruction_decode/add_358/carry [3]), .CO(
        \instruction_decode/add_358/carry [4]), .S(\instruction_decode/N11 )
         );
  ADD32 \instruction_decode/add_358/U1_4  ( .A(pc_out[4]), .B(inst_out[2]), 
        .CI(\instruction_decode/add_358/carry [4]), .CO(
        \instruction_decode/add_358/carry [5]), .S(\instruction_decode/N12 )
         );
  ADD32 \instruction_decode/add_358/U1_5  ( .A(pc_out[5]), .B(inst_out[3]), 
        .CI(\instruction_decode/add_358/carry [5]), .CO(
        \instruction_decode/add_358/carry [6]), .S(\instruction_decode/N13 )
         );
  ADD32 \instruction_decode/add_358/U1_6  ( .A(pc_out[6]), .B(inst_out[4]), 
        .CI(\instruction_decode/add_358/carry [6]), .CO(
        \instruction_decode/add_358/carry [7]), .S(\instruction_decode/N14 )
         );
  ADD32 \instruction_decode/add_358/U1_7  ( .A(pc_out[7]), .B(inst_out[5]), 
        .CI(\instruction_decode/add_358/carry [7]), .CO(
        \instruction_decode/add_358/carry [8]), .S(\instruction_decode/N15 )
         );
  ADD32 \instruction_decode/add_358/U1_8  ( .A(pc_out[8]), .B(inst_out[6]), 
        .CI(\instruction_decode/add_358/carry [8]), .CO(
        \instruction_decode/add_358/carry [9]), .S(\instruction_decode/N16 )
         );
  ADD32 \instruction_decode/add_358/U1_9  ( .A(pc_out[9]), .B(inst_out[7]), 
        .CI(\instruction_decode/add_358/carry [9]), .CO(
        \instruction_decode/add_358/carry [10]), .S(\instruction_decode/N17 )
         );
  ADD32 \instruction_decode/add_358/U1_10  ( .A(pc_out[10]), .B(inst_out[8]), 
        .CI(\instruction_decode/add_358/carry [10]), .CO(
        \instruction_decode/add_358/carry [11]), .S(\instruction_decode/N18 )
         );
  ADD32 \instruction_decode/add_358/U1_11  ( .A(pc_out[11]), .B(inst_out[9]), 
        .CI(\instruction_decode/add_358/carry [11]), .CO(
        \instruction_decode/add_358/carry [12]), .S(\instruction_decode/N19 )
         );
  ADD32 \instruction_decode/add_358/U1_12  ( .A(pc_out[12]), .B(inst_out[10]), 
        .CI(\instruction_decode/add_358/carry [12]), .CO(
        \instruction_decode/add_358/carry [13]), .S(\instruction_decode/N20 )
         );
  ADD32 \instruction_decode/add_358/U1_13  ( .A(pc_out[13]), .B(inst_out[11]), 
        .CI(\instruction_decode/add_358/carry [13]), .CO(
        \instruction_decode/add_358/carry [14]), .S(\instruction_decode/N21 )
         );
  ADD32 \instruction_decode/add_358/U1_14  ( .A(pc_out[14]), .B(inst_out[12]), 
        .CI(\instruction_decode/add_358/carry [14]), .CO(
        \instruction_decode/add_358/carry [15]), .S(\instruction_decode/N22 )
         );
  DF3 \execute/write_data_ex_reg[0]  ( .D(\execute/op_21 [0]), .C(clk), .Q(
        ram_data[0]) );
  DF3 \execute/write_data_ex_reg[1]  ( .D(\execute/op_21 [1]), .C(clk), .Q(
        ram_data[1]) );
  DF3 \execute/write_data_ex_reg[2]  ( .D(\execute/op_21 [2]), .C(clk), .Q(
        ram_data[2]) );
  DF3 \execute/write_data_ex_reg[3]  ( .D(n5813), .C(clk), .Q(ram_data[3]) );
  DF3 \execute/write_data_ex_reg[4]  ( .D(\execute/op_21 [4]), .C(clk), .Q(
        ram_data[4]) );
  DF3 \execute/write_data_ex_reg[5]  ( .D(\execute/op_21 [5]), .C(clk), .Q(
        ram_data[5]) );
  DF3 \execute/write_data_ex_reg[6]  ( .D(\execute/op_21 [6]), .C(clk), .Q(
        ram_data[6]) );
  DF3 \execute/write_data_ex_reg[7]  ( .D(\execute/op_21 [7]), .C(clk), .Q(
        ram_data[7]) );
  DF3 \execute/write_data_ex_reg[8]  ( .D(\execute/op_21 [8]), .C(clk), .Q(
        ram_data[8]) );
  DF3 \execute/write_data_ex_reg[9]  ( .D(\execute/op_21 [9]), .C(clk), .Q(
        ram_data[9]) );
  DF3 \execute/write_data_ex_reg[10]  ( .D(\execute/op_21 [10]), .C(clk), .Q(
        ram_data[10]) );
  DF3 \execute/write_data_ex_reg[11]  ( .D(\execute/op_21 [11]), .C(clk), .Q(
        ram_data[11]) );
  DF3 \execute/write_data_ex_reg[12]  ( .D(\execute/op_21 [12]), .C(clk), .Q(
        ram_data[12]) );
  DF3 \execute/write_data_ex_reg[13]  ( .D(\execute/op_21 [13]), .C(clk), .Q(
        ram_data[13]) );
  DF3 \execute/write_data_ex_reg[14]  ( .D(\execute/op_21 [14]), .C(clk), .Q(
        ram_data[14]) );
  DF3 \execute/write_data_ex_reg[15]  ( .D(\execute/op_21 [15]), .C(clk), .Q(
        ram_data[15]) );
  DF3 \execute/write_data_ex_reg[16]  ( .D(\execute/op_21 [16]), .C(clk), .Q(
        ram_data[16]) );
  DF3 \execute/write_data_ex_reg[17]  ( .D(\execute/op_21 [17]), .C(clk), .Q(
        ram_data[17]) );
  DF3 \execute/write_data_ex_reg[18]  ( .D(\execute/op_21 [18]), .C(clk), .Q(
        ram_data[18]) );
  DF3 \execute/write_data_ex_reg[19]  ( .D(\execute/op_21 [19]), .C(clk), .Q(
        ram_data[19]) );
  DF3 \execute/write_data_ex_reg[20]  ( .D(\execute/op_21 [20]), .C(clk), .Q(
        ram_data[20]) );
  DF3 \execute/write_data_ex_reg[21]  ( .D(\execute/op_21 [21]), .C(clk), .Q(
        ram_data[21]) );
  DF3 \execute/write_data_ex_reg[22]  ( .D(\execute/op_21 [22]), .C(clk), .Q(
        ram_data[22]) );
  DF3 \execute/write_data_ex_reg[23]  ( .D(\execute/op_21 [23]), .C(clk), .Q(
        ram_data[23]) );
  DF3 \execute/write_data_ex_reg[24]  ( .D(\execute/op_21 [24]), .C(clk), .Q(
        ram_data[24]) );
  DF3 \execute/write_data_ex_reg[25]  ( .D(\execute/op_21 [25]), .C(clk), .Q(
        ram_data[25]) );
  DF3 \execute/write_data_ex_reg[26]  ( .D(\execute/op_21 [26]), .C(clk), .Q(
        ram_data[26]) );
  DF3 \execute/write_data_ex_reg[27]  ( .D(\execute/op_21 [27]), .C(clk), .Q(
        ram_data[27]) );
  DF3 \execute/write_data_ex_reg[28]  ( .D(\execute/op_21 [28]), .C(clk), .Q(
        ram_data[28]) );
  DF3 \execute/write_data_ex_reg[29]  ( .D(\execute/op_21 [29]), .C(clk), .Q(
        ram_data[29]) );
  DF3 \execute/write_data_ex_reg[30]  ( .D(\execute/op_21 [30]), .C(clk), .Q(
        ram_data[30]) );
  DF3 \execute/write_data_ex_reg[31]  ( .D(\execute/op_21 [31]), .C(clk), .Q(
        ram_data[31]) );
  DF3 \execute/res_reg[31]  ( .D(\execute/old_res [31]), .C(clk), .Q(
        ram_adr[31]) );
  DF3 \execute/res_reg[30]  ( .D(\execute/old_res [30]), .C(clk), .Q(
        ram_adr[30]) );
  DF3 \execute/res_reg[29]  ( .D(\execute/old_res [29]), .C(clk), .Q(
        ram_adr[29]) );
  DF3 \execute/res_reg[28]  ( .D(\execute/old_res [28]), .C(clk), .Q(
        ram_adr[28]) );
  DF3 \execute/res_reg[27]  ( .D(\execute/old_res [27]), .C(clk), .Q(
        ram_adr[27]) );
  DF3 \execute/res_reg[26]  ( .D(\execute/old_res [26]), .C(clk), .Q(
        ram_adr[26]) );
  DF3 \execute/res_reg[25]  ( .D(\execute/old_res [25]), .C(clk), .Q(
        ram_adr[25]) );
  DF3 \execute/res_reg[24]  ( .D(\execute/old_res [24]), .C(clk), .Q(
        ram_adr[24]) );
  DF3 \execute/res_reg[23]  ( .D(\execute/old_res [23]), .C(clk), .Q(
        ram_adr[23]) );
  DF3 \execute/res_reg[22]  ( .D(n1220), .C(clk), .Q(ram_adr[22]) );
  DF3 \execute/res_reg[21]  ( .D(\execute/old_res [21]), .C(clk), .Q(
        ram_adr[21]) );
  DF3 \execute/res_reg[20]  ( .D(\execute/old_res [20]), .C(clk), .Q(
        ram_adr[20]) );
  DF3 \execute/res_reg[19]  ( .D(\execute/old_res [19]), .C(clk), .Q(
        ram_adr[19]) );
  DF3 \execute/res_reg[18]  ( .D(n1217), .C(clk), .Q(ram_adr[18]) );
  DF3 \execute/res_reg[17]  ( .D(\execute/old_res [17]), .C(clk), .Q(
        ram_adr[17]) );
  DF3 \execute/res_reg[16]  ( .D(\execute/old_res [16]), .C(clk), .Q(
        ram_adr[16]) );
  DF3 \execute/res_reg[15]  ( .D(\execute/old_res [15]), .C(clk), .Q(
        ram_adr[15]) );
  DF3 \execute/res_reg[14]  ( .D(\execute/old_res [14]), .C(clk), .Q(
        ram_adr[14]) );
  DF3 \execute/res_reg[13]  ( .D(\execute/old_res [13]), .C(clk), .Q(
        ram_adr[13]) );
  DF3 \execute/res_reg[12]  ( .D(\execute/old_res [12]), .C(clk), .Q(
        ram_adr[12]) );
  DF3 \execute/res_reg[11]  ( .D(\execute/old_res [11]), .C(clk), .Q(
        ram_adr[11]) );
  DF3 \execute/res_reg[10]  ( .D(\execute/old_res [10]), .C(clk), .Q(
        ram_adr[10]) );
  DF3 \execute/res_reg[9]  ( .D(\execute/old_res [9]), .C(clk), .Q(ram_adr[9])
         );
  DF3 \execute/res_reg[8]  ( .D(\execute/old_res [8]), .C(clk), .Q(ram_adr[8])
         );
  DF3 \execute/res_reg[7]  ( .D(\execute/old_res [7]), .C(clk), .Q(ram_adr[7])
         );
  DF3 \execute/res_reg[6]  ( .D(\execute/old_res [6]), .C(clk), .Q(ram_adr[6])
         );
  DF3 \execute/res_reg[5]  ( .D(\execute/old_res [5]), .C(clk), .Q(ram_adr[5])
         );
  DF3 \execute/res_reg[4]  ( .D(\execute/old_res [4]), .C(clk), .Q(ram_adr[4])
         );
  DF3 \execute/res_reg[3]  ( .D(\execute/old_res [3]), .C(clk), .Q(ram_adr[3])
         );
  DF3 \execute/res_reg[2]  ( .D(\execute/old_res [2]), .C(clk), .Q(ram_adr[2])
         );
  DF3 \execute/res_reg[1]  ( .D(\execute/old_res [1]), .C(clk), .Q(ram_adr[1])
         );
  DF3 \execute/res_reg[0]  ( .D(\execute/old_res [0]), .C(clk), .Q(ram_adr[0])
         );
  DF3 \execute/write_register_ex_reg[0]  ( .D(n5803), .C(clk), .Q(
        write_register_ex[0]) );
  DF3 \execute/write_register_ex_reg[1]  ( .D(n5804), .C(clk), .Q(
        write_register_ex[1]) );
  DF3 \execute/write_register_ex_reg[2]  ( .D(n5805), .C(clk), .Q(
        write_register_ex[2]), .QN(n6227) );
  DF3 \execute/write_register_ex_reg[3]  ( .D(n5806), .C(clk), .Q(
        write_register_ex[3]), .QN(n6226) );
  DF3 \execute/write_register_ex_reg[4]  ( .D(n5807), .C(clk), .Q(
        write_register_ex[4]), .QN(n6268) );
  DF3 \execute/wb_MEM_reg[0]  ( .D(n5768), .C(clk), .Q(wb_MEM[0]) );
  DF3 \execute/wb_MEM_reg[1]  ( .D(n5767), .C(clk), .Q(wb_MEM[1]) );
  DF3 \execute/m_MEM_reg[0]  ( .D(n5769), .C(clk), .Q(ram_write) );
  DF3 \execute/m_MEM_reg[1]  ( .D(n5770), .C(clk), .Q(ram_read) );
  DF3 \execute/m_MEM_reg[2]  ( .D(n5771), .C(clk), .Q(ram_size[0]) );
  DF3 \execute/m_MEM_reg[3]  ( .D(n5772), .C(clk), .Q(ram_size[1]) );
  DF3 \memory/read_data_reg[0]  ( .D(ram_word[0]), .C(clk), .QN(n5658) );
  DF3 \memory/address_WB_reg[0]  ( .D(ram_adr[0]), .C(clk), .QN(n5659) );
  DF3 \memory/address_WB_reg[4]  ( .D(ram_adr[4]), .C(clk), .QN(n5645) );
  DF3 \memory/write_register_mem_reg[0]  ( .D(write_register_ex[0]), .C(clk), 
        .Q(write_register[0]), .QN(n5867) );
  DF3 \memory/write_register_mem_reg[1]  ( .D(write_register_ex[1]), .C(clk), 
        .Q(write_register[1]), .QN(n5848) );
  DF3 \memory/write_register_mem_reg[2]  ( .D(write_register_ex[2]), .C(clk), 
        .Q(write_register[2]), .QN(n5941) );
  DF3 \memory/write_register_mem_reg[3]  ( .D(write_register_ex[3]), .C(clk), 
        .Q(write_register[3]), .QN(n6069) );
  DF3 \memory/write_register_mem_reg[4]  ( .D(write_register_ex[4]), .C(clk), 
        .Q(write_register[4]), .QN(n5943) );
  DF3 \memory/wb_reg[0]  ( .D(wb_MEM[0]), .C(clk), .Q(\wb_WB[0] ), .QN(n6068)
         );
  DF3 \memory/wb_reg[1]  ( .D(wb_MEM[1]), .C(clk), .Q(reg_write) );
  OAI212 U42 ( .A(n5716), .B(n5945), .C(n6279), .Q(n1769) );
  OAI212 U43 ( .A(n6286), .B(n1774), .C(n1775), .Q(n5774) );
  OAI212 U61 ( .A(n5826), .B(n1156), .C(n1794), .Q(n5780) );
  OAI212 U68 ( .A(n6288), .B(n1800), .C(n1801), .Q(n5783) );
  OAI212 U71 ( .A(n6288), .B(n1803), .C(n1804), .Q(n5784) );
  OAI212 U74 ( .A(n6300), .B(n1806), .C(n1807), .Q(n5785) );
  OAI212 U77 ( .A(n6287), .B(n1809), .C(n1810), .Q(n5786) );
  OAI212 U80 ( .A(n6286), .B(n1812), .C(n1813), .Q(n5787) );
  OAI212 U87 ( .A(n6291), .B(n1817), .C(n1818), .Q(n5790) );
  OAI212 U90 ( .A(n6292), .B(n1820), .C(n1821), .Q(n5791) );
  OAI212 U105 ( .A(n6298), .B(n1835), .C(n1836), .Q(n5796) );
  OAI212 U108 ( .A(n6299), .B(\instruction_fetch/n87 ), .C(n1838), .Q(n5797)
         );
  OAI212 U112 ( .A(n6274), .B(n1842), .C(n1843), .Q(n5798) );
  OAI212 U115 ( .A(n6294), .B(n1845), .C(n1846), .Q(n5799) );
  OAI222 U118 ( .A(n6313), .B(n4575), .C(n6301), .D(n1848), .Q(n5800) );
  OAI222 U124 ( .A(n1465), .B(n5626), .C(n1485), .D(n1854), .Q(n5803) );
  OAI222 U125 ( .A(n1465), .B(n5625), .C(n6209), .D(n1854), .Q(n5804) );
  OAI222 U126 ( .A(n1465), .B(n5624), .C(n6091), .D(n1854), .Q(n5805) );
  OAI222 U127 ( .A(n1465), .B(n5623), .C(n1489), .D(n1854), .Q(n5806) );
  OAI222 U128 ( .A(n1465), .B(n5622), .C(n1490), .D(n1854), .Q(n5807) );
  OAI212 U130 ( .A(n6292), .B(n1857), .C(n1858), .Q(
        \instruction_fetch/pc_4 [8]) );
  OAI2112 U167 ( .A(n1865), .B(n1185), .C(n1147), .D(n1866), .Q(n1780) );
  AOI222 U168 ( .A(\instruction_decode/old_ex [2]), .B(n1160), .C(n1868), .D(
        \instruction_decode/old_ex [1]), .Q(n1867) );
  OAI222 U214 ( .A(n1919), .B(n6499), .C(n6320), .D(n1920), .Q(n1918) );
  OAI222 U216 ( .A(n4907), .B(n6590), .C(n4906), .D(n6582), .Q(n1924) );
  OAI222 U217 ( .A(n5151), .B(n6580), .C(n5150), .D(n1928), .Q(n1923) );
  OAI222 U218 ( .A(n5153), .B(n6565), .C(n5152), .D(n6564), .Q(n1922) );
  OAI222 U219 ( .A(n5155), .B(n6556), .C(n5154), .D(n1932), .Q(n1921) );
  OAI222 U221 ( .A(n4857), .B(n6590), .C(n4856), .D(n6583), .Q(n1936) );
  OAI222 U225 ( .A(n4693), .B(n6419), .C(n4692), .D(n6421), .Q(n1917) );
  OAI212 U227 ( .A(n6402), .B(n5972), .C(n1942), .Q(n1915) );
  OAI222 U230 ( .A(n1170), .B(n6018), .C(n6401), .D(n5897), .Q(n1947) );
  OAI222 U231 ( .A(n4746), .B(n6393), .C(n6399), .D(n5998), .Q(n1946) );
  OAI222 U293 ( .A(n1978), .B(n1974), .C(n1979), .D(n1972), .Q(
        \instruction_decode/old_ex [2]) );
  OAI212 U304 ( .A(n1975), .B(n1984), .C(n1970), .Q(n1967) );
  OAI312 U309 ( .A(n1145), .B(n5730), .C(n1187), .D(n1973), .Q(n1983) );
  AOI2112 U315 ( .A(n6280), .B(n1413), .C(n1988), .D(n5700), .Q(n1987) );
  AOI312 U316 ( .A(n1989), .B(n1461), .C(n6280), .D(n1990), .Q(n1988) );
  OAI222 U321 ( .A(n2002), .B(n6493), .C(n6317), .D(n2003), .Q(n2001) );
  OAI222 U323 ( .A(n5319), .B(n6548), .C(n5318), .D(n6546), .Q(n2007) );
  OAI222 U324 ( .A(n5201), .B(n6539), .C(n5200), .D(n6537), .Q(n2006) );
  OAI222 U325 ( .A(n5203), .B(n6530), .C(n5202), .D(n6527), .Q(n2005) );
  OAI222 U326 ( .A(n5205), .B(n6526), .C(n5204), .D(n6518), .Q(n2004) );
  OAI222 U328 ( .A(n4873), .B(n6553), .C(n4872), .D(n6546), .Q(n2019) );
  OAI222 U329 ( .A(n5047), .B(n6544), .C(n5046), .D(n6537), .Q(n2018) );
  OAI222 U331 ( .A(n5341), .B(n6526), .C(n5340), .D(n6518), .Q(n2016) );
  OAI222 U332 ( .A(n4633), .B(n6483), .C(n4632), .D(n6485), .Q(n2000) );
  OAI222 U333 ( .A(n4631), .B(n6479), .C(n4630), .D(n6481), .Q(n1999) );
  OAI212 U334 ( .A(n6467), .B(n5971), .C(n2025), .Q(n1998) );
  OAI222 U337 ( .A(n1162), .B(n6017), .C(n6462), .D(n5857), .Q(n2030) );
  OAI222 U338 ( .A(n4774), .B(n6456), .C(n6458), .D(n5997), .Q(n2029) );
  OAI222 U343 ( .A(n2046), .B(n6493), .C(n6318), .D(n2047), .Q(n2045) );
  OAI222 U350 ( .A(n4897), .B(n6553), .C(n4896), .D(n6546), .Q(n2055) );
  OAI222 U354 ( .A(n4637), .B(n6482), .C(n4636), .D(n6484), .Q(n2044) );
  OAI222 U355 ( .A(n4635), .B(n6478), .C(n4634), .D(n6480), .Q(n2043) );
  OAI212 U356 ( .A(n6466), .B(n5970), .C(n2056), .Q(n2042) );
  OAI222 U359 ( .A(n1162), .B(n6016), .C(n6464), .D(n5896), .Q(n2058) );
  OAI222 U360 ( .A(n4806), .B(n6455), .C(n6457), .D(n5996), .Q(n2057) );
  OAI222 U365 ( .A(n2067), .B(n6493), .C(n6316), .D(n2068), .Q(n2066) );
  OAI222 U372 ( .A(n4917), .B(n6553), .C(n4916), .D(n6546), .Q(n2076) );
  OAI222 U376 ( .A(n4641), .B(n2020), .C(n4640), .D(n2021), .Q(n2065) );
  OAI212 U378 ( .A(n2024), .B(n5969), .C(n2077), .Q(n2063) );
  OAI222 U381 ( .A(n1162), .B(n6015), .C(n6464), .D(n5895), .Q(n2079) );
  OAI222 U382 ( .A(n4822), .B(n2032), .C(n2033), .D(n5995), .Q(n2078) );
  OAI222 U387 ( .A(n2088), .B(n6493), .C(n6316), .D(n2089), .Q(n2087) );
  OAI222 U389 ( .A(n4919), .B(n6553), .C(n4918), .D(n6546), .Q(n2093) );
  OAI222 U390 ( .A(n5189), .B(n6544), .C(n5188), .D(n6537), .Q(n2092) );
  OAI222 U391 ( .A(n5191), .B(n6535), .C(n5190), .D(n2013), .Q(n2091) );
  OAI222 U392 ( .A(n5193), .B(n6526), .C(n5192), .D(n2015), .Q(n2090) );
  OAI222 U394 ( .A(n4867), .B(n6553), .C(n4866), .D(n6546), .Q(n2097) );
  OAI222 U395 ( .A(n5029), .B(n6544), .C(n5028), .D(n6537), .Q(n2096) );
  OAI222 U396 ( .A(n5031), .B(n6535), .C(n5030), .D(n2013), .Q(n2095) );
  OAI222 U397 ( .A(n5033), .B(n6526), .C(n5032), .D(n6519), .Q(n2094) );
  OAI222 U398 ( .A(n4645), .B(n6483), .C(n4644), .D(n6485), .Q(n2086) );
  OAI222 U399 ( .A(n4643), .B(n6479), .C(n4642), .D(n6481), .Q(n2085) );
  OAI212 U400 ( .A(n6467), .B(n5968), .C(n2098), .Q(n2084) );
  OAI222 U403 ( .A(n1162), .B(n6014), .C(n6463), .D(n5894), .Q(n2100) );
  OAI222 U404 ( .A(n4766), .B(n6456), .C(n6458), .D(n5994), .Q(n2099) );
  OAI222 U409 ( .A(n2109), .B(n6493), .C(n6316), .D(n2110), .Q(n2108) );
  OAI222 U411 ( .A(n4933), .B(n6553), .C(n4932), .D(n6546), .Q(n2114) );
  OAI222 U412 ( .A(n5235), .B(n6544), .C(n5234), .D(n6537), .Q(n2113) );
  OAI222 U413 ( .A(n5237), .B(n6535), .C(n5236), .D(n2013), .Q(n2112) );
  OAI222 U414 ( .A(n5239), .B(n6526), .C(n5238), .D(n2015), .Q(n2111) );
  OAI222 U416 ( .A(n4887), .B(n6553), .C(n4886), .D(n6546), .Q(n2118) );
  OAI222 U417 ( .A(n5087), .B(n6544), .C(n5086), .D(n6537), .Q(n2117) );
  OAI222 U418 ( .A(n5089), .B(n6535), .C(n5088), .D(n2013), .Q(n2116) );
  OAI222 U419 ( .A(n5091), .B(n6526), .C(n5090), .D(n6518), .Q(n2115) );
  OAI222 U420 ( .A(n4649), .B(n6482), .C(n4648), .D(n6484), .Q(n2107) );
  OAI222 U421 ( .A(n4647), .B(n6478), .C(n4646), .D(n6480), .Q(n2106) );
  OAI212 U422 ( .A(n6466), .B(n5967), .C(n2119), .Q(n2105) );
  OAI222 U425 ( .A(n1162), .B(n6013), .C(n6463), .D(n5893), .Q(n2121) );
  OAI222 U426 ( .A(n4794), .B(n6455), .C(n6457), .D(n5993), .Q(n2120) );
  OAI222 U431 ( .A(n2130), .B(n6493), .C(n6316), .D(n2131), .Q(n2129) );
  OAI222 U433 ( .A(n4945), .B(n6552), .C(n4944), .D(n6546), .Q(n2135) );
  OAI222 U434 ( .A(n5271), .B(n6543), .C(n5270), .D(n6537), .Q(n2134) );
  OAI222 U435 ( .A(n5273), .B(n6534), .C(n5272), .D(n6528), .Q(n2133) );
  OAI222 U436 ( .A(n5345), .B(n6525), .C(n5344), .D(n6519), .Q(n2132) );
  OAI222 U438 ( .A(n4909), .B(n6552), .C(n4908), .D(n6546), .Q(n2139) );
  OAI222 U439 ( .A(n5157), .B(n6543), .C(n5156), .D(n6537), .Q(n2138) );
  OAI222 U441 ( .A(n5327), .B(n6525), .C(n5326), .D(n6519), .Q(n2136) );
  OAI222 U442 ( .A(n4653), .B(n2020), .C(n4652), .D(n2021), .Q(n2128) );
  OAI222 U443 ( .A(n4651), .B(n2022), .C(n4650), .D(n2023), .Q(n2127) );
  OAI212 U444 ( .A(n2024), .B(n5966), .C(n2140), .Q(n2126) );
  OAI222 U447 ( .A(n1162), .B(n6012), .C(n6460), .D(n5892), .Q(n2142) );
  OAI222 U448 ( .A(n4818), .B(n2032), .C(n2033), .D(n5992), .Q(n2141) );
  OAI222 U453 ( .A(n2151), .B(n6493), .C(n6318), .D(n2152), .Q(n2150) );
  OAI222 U455 ( .A(n5321), .B(n6552), .C(n5320), .D(n2009), .Q(n2156) );
  OAI222 U456 ( .A(n5281), .B(n6543), .C(n5280), .D(n2011), .Q(n2155) );
  OAI222 U457 ( .A(n5283), .B(n6534), .C(n5282), .D(n2013), .Q(n2154) );
  OAI222 U458 ( .A(n5285), .B(n6525), .C(n5284), .D(n2015), .Q(n2153) );
  OAI222 U460 ( .A(n4925), .B(n6552), .C(n4924), .D(n2009), .Q(n2160) );
  OAI222 U461 ( .A(n5213), .B(n6543), .C(n5212), .D(n2011), .Q(n2159) );
  OAI222 U462 ( .A(n5215), .B(n6534), .C(n5214), .D(n2013), .Q(n2158) );
  OAI222 U463 ( .A(n5317), .B(n6525), .C(n5316), .D(n2015), .Q(n2157) );
  OAI222 U464 ( .A(n4657), .B(n6483), .C(n4656), .D(n6485), .Q(n2149) );
  OAI222 U465 ( .A(n4655), .B(n6479), .C(n4654), .D(n6481), .Q(n2148) );
  OAI212 U466 ( .A(n6467), .B(n5965), .C(n2161), .Q(n2147) );
  OAI222 U469 ( .A(n1162), .B(n6011), .C(n6462), .D(n5891), .Q(n2163) );
  OAI222 U470 ( .A(n4826), .B(n6456), .C(n6458), .D(n5991), .Q(n2162) );
  OAI222 U475 ( .A(n2172), .B(n6493), .C(n6316), .D(n2173), .Q(n2171) );
  OAI222 U477 ( .A(n4935), .B(n6552), .C(n4934), .D(n2009), .Q(n2177) );
  OAI222 U478 ( .A(n5241), .B(n6543), .C(n5240), .D(n2011), .Q(n2176) );
  OAI222 U479 ( .A(n5243), .B(n6534), .C(n5242), .D(n2013), .Q(n2175) );
  OAI222 U480 ( .A(n5245), .B(n6525), .C(n5244), .D(n2015), .Q(n2174) );
  OAI222 U482 ( .A(n4889), .B(n6552), .C(n4888), .D(n2009), .Q(n2181) );
  OAI222 U483 ( .A(n5099), .B(n6543), .C(n5098), .D(n2011), .Q(n2180) );
  OAI222 U484 ( .A(n5101), .B(n6534), .C(n5100), .D(n2013), .Q(n2179) );
  OAI222 U485 ( .A(n5103), .B(n6525), .C(n5102), .D(n2015), .Q(n2178) );
  OAI222 U486 ( .A(n4585), .B(n6482), .C(n4584), .D(n6484), .Q(n2170) );
  OAI222 U487 ( .A(n4583), .B(n6478), .C(n4582), .D(n6480), .Q(n2169) );
  OAI212 U488 ( .A(n6466), .B(n5873), .C(n2182), .Q(n2168) );
  OAI222 U491 ( .A(n1162), .B(n5939), .C(n2031), .D(n5858), .Q(n2184) );
  OAI222 U492 ( .A(n4798), .B(n6455), .C(n6457), .D(n5890), .Q(n2183) );
  OAI222 U497 ( .A(n2193), .B(n6493), .C(n6316), .D(n2194), .Q(n2192) );
  OAI222 U499 ( .A(n4853), .B(n6552), .C(n4852), .D(n6545), .Q(n2198) );
  OAI222 U500 ( .A(n4991), .B(n6543), .C(n4990), .D(n6537), .Q(n2197) );
  OAI222 U501 ( .A(n4993), .B(n6534), .C(n4992), .D(n2013), .Q(n2196) );
  OAI222 U502 ( .A(n4995), .B(n6525), .C(n4994), .D(n6518), .Q(n2195) );
  OAI222 U504 ( .A(n4839), .B(n6552), .C(n4838), .D(n2009), .Q(n2202) );
  OAI222 U505 ( .A(n4953), .B(n6543), .C(n4952), .D(n2011), .Q(n2201) );
  OAI222 U506 ( .A(n4955), .B(n6534), .C(n4954), .D(n2013), .Q(n2200) );
  OAI222 U507 ( .A(n4957), .B(n6525), .C(n4956), .D(n2015), .Q(n2199) );
  OAI222 U508 ( .A(n4589), .B(n2020), .C(n4588), .D(n2021), .Q(n2191) );
  OAI212 U510 ( .A(n2024), .B(n5964), .C(n2203), .Q(n2189) );
  OAI222 U514 ( .A(n4710), .B(n2032), .C(n2033), .D(n5990), .Q(n2204) );
  OAI222 U519 ( .A(n2214), .B(n6494), .C(n6316), .D(n2215), .Q(n2213) );
  OAI222 U521 ( .A(n4921), .B(n6552), .C(n4920), .D(n2009), .Q(n2219) );
  OAI222 U522 ( .A(n5195), .B(n6543), .C(n5194), .D(n2011), .Q(n2218) );
  OAI222 U523 ( .A(n5197), .B(n6534), .C(n5196), .D(n2013), .Q(n2217) );
  OAI222 U524 ( .A(n5199), .B(n6525), .C(n5198), .D(n2015), .Q(n2216) );
  OAI222 U527 ( .A(n5035), .B(n6542), .C(n5034), .D(n2011), .Q(n2222) );
  OAI222 U528 ( .A(n5037), .B(n6533), .C(n5036), .D(n2013), .Q(n2221) );
  OAI222 U529 ( .A(n5039), .B(n6524), .C(n5038), .D(n2015), .Q(n2220) );
  OAI222 U530 ( .A(n4661), .B(n6483), .C(n4660), .D(n6485), .Q(n2212) );
  OAI222 U531 ( .A(n4659), .B(n6479), .C(n4658), .D(n6481), .Q(n2211) );
  OAI212 U532 ( .A(n6467), .B(n5963), .C(n2224), .Q(n2210) );
  OAI222 U535 ( .A(n1162), .B(n6066), .C(n6464), .D(n5840), .Q(n2226) );
  OAI222 U536 ( .A(n4770), .B(n6456), .C(n6458), .D(n5989), .Q(n2225) );
  OAI222 U541 ( .A(n2235), .B(n6493), .C(n6316), .D(n2236), .Q(n2234) );
  OAI222 U543 ( .A(n4871), .B(n6551), .C(n4870), .D(n6546), .Q(n2240) );
  OAI222 U544 ( .A(n5041), .B(n6542), .C(n5040), .D(n6536), .Q(n2239) );
  OAI222 U545 ( .A(n5043), .B(n6533), .C(n5042), .D(n6528), .Q(n2238) );
  OAI222 U546 ( .A(n5045), .B(n6524), .C(n5044), .D(n6519), .Q(n2237) );
  OAI222 U548 ( .A(n4841), .B(n6551), .C(n4840), .D(n2009), .Q(n2244) );
  OAI222 U549 ( .A(n4959), .B(n6542), .C(n4958), .D(n2011), .Q(n2243) );
  OAI222 U550 ( .A(n4961), .B(n6533), .C(n4960), .D(n2013), .Q(n2242) );
  OAI222 U552 ( .A(n4593), .B(n6482), .C(n4592), .D(n6484), .Q(n2233) );
  OAI222 U553 ( .A(n4591), .B(n6478), .C(n4590), .D(n6480), .Q(n2232) );
  OAI212 U554 ( .A(n6466), .B(n5962), .C(n2245), .Q(n2231) );
  OAI222 U557 ( .A(n1162), .B(n6065), .C(n6464), .D(n5907), .Q(n2247) );
  OAI222 U558 ( .A(n4714), .B(n6455), .C(n6457), .D(n5988), .Q(n2246) );
  OAI222 U563 ( .A(n2256), .B(n6493), .C(n6316), .D(n2257), .Q(n2255) );
  OAI222 U565 ( .A(n4895), .B(n6551), .C(n4894), .D(n2009), .Q(n2261) );
  OAI222 U566 ( .A(n5117), .B(n6542), .C(n5116), .D(n2011), .Q(n2260) );
  OAI222 U567 ( .A(n5119), .B(n6533), .C(n5118), .D(n2013), .Q(n2259) );
  OAI222 U568 ( .A(n5121), .B(n6524), .C(n5120), .D(n2015), .Q(n2258) );
  OAI222 U570 ( .A(n4849), .B(n6551), .C(n4848), .D(n2009), .Q(n2265) );
  OAI222 U571 ( .A(n4983), .B(n6542), .C(n4982), .D(n2011), .Q(n2264) );
  OAI222 U572 ( .A(n4985), .B(n6533), .C(n4984), .D(n2013), .Q(n2263) );
  OAI222 U573 ( .A(n5351), .B(n6524), .C(n5350), .D(n2015), .Q(n2262) );
  OAI222 U574 ( .A(n4597), .B(n2020), .C(n4596), .D(n2021), .Q(n2254) );
  OAI222 U575 ( .A(n4595), .B(n2022), .C(n4594), .D(n2023), .Q(n2253) );
  OAI212 U576 ( .A(n2024), .B(n5961), .C(n2266), .Q(n2252) );
  OAI222 U579 ( .A(n1162), .B(n6064), .C(n6463), .D(n5906), .Q(n2268) );
  OAI222 U580 ( .A(n4734), .B(n2032), .C(n2033), .D(n5987), .Q(n2267) );
  OAI222 U585 ( .A(n2277), .B(n6494), .C(n6316), .D(n2278), .Q(n2276) );
  OAI222 U587 ( .A(n4915), .B(n6551), .C(n4914), .D(n2009), .Q(n2282) );
  OAI222 U588 ( .A(n5173), .B(n6542), .C(n5172), .D(n2011), .Q(n2281) );
  OAI222 U589 ( .A(n5175), .B(n6533), .C(n5174), .D(n2013), .Q(n2280) );
  OAI222 U590 ( .A(n5335), .B(n6524), .C(n5334), .D(n2015), .Q(n2279) );
  OAI222 U592 ( .A(n4863), .B(n6551), .C(n4862), .D(n6545), .Q(n2286) );
  OAI222 U593 ( .A(n5017), .B(n6542), .C(n5016), .D(n2011), .Q(n2285) );
  OAI222 U594 ( .A(n5019), .B(n6533), .C(n5018), .D(n6528), .Q(n2284) );
  OAI222 U595 ( .A(n5021), .B(n6524), .C(n5020), .D(n6518), .Q(n2283) );
  OAI222 U596 ( .A(n4601), .B(n6483), .C(n4600), .D(n6485), .Q(n2275) );
  OAI222 U597 ( .A(n4599), .B(n6479), .C(n4598), .D(n6481), .Q(n2274) );
  OAI212 U598 ( .A(n6467), .B(n5960), .C(n2287), .Q(n2273) );
  OAI222 U601 ( .A(n1162), .B(n6010), .C(n6460), .D(n5889), .Q(n2289) );
  OAI222 U602 ( .A(n4758), .B(n6456), .C(n6458), .D(n5986), .Q(n2288) );
  OAI222 U607 ( .A(n2298), .B(n6494), .C(n6316), .D(n2299), .Q(n2297) );
  OAI222 U612 ( .A(n5061), .B(n6524), .C(n5060), .D(n2015), .Q(n2300) );
  OAI222 U614 ( .A(n4843), .B(n6551), .C(n4842), .D(n2009), .Q(n2307) );
  OAI222 U618 ( .A(n4605), .B(n6482), .C(n4604), .D(n6484), .Q(n2296) );
  OAI212 U620 ( .A(n6466), .B(n5959), .C(n2308), .Q(n2294) );
  OAI222 U623 ( .A(n1162), .B(n6063), .C(n6460), .D(n5905), .Q(n2310) );
  OAI222 U624 ( .A(n4718), .B(n6455), .C(n6457), .D(n5985), .Q(n2309) );
  OAI222 U629 ( .A(n2319), .B(n6494), .C(n6316), .D(n2320), .Q(n2318) );
  OAI222 U631 ( .A(n4899), .B(n6550), .C(n4898), .D(n6545), .Q(n2324) );
  OAI222 U632 ( .A(n5129), .B(n6541), .C(n5128), .D(n6537), .Q(n2323) );
  OAI222 U633 ( .A(n5131), .B(n6532), .C(n5130), .D(n6528), .Q(n2322) );
  OAI222 U634 ( .A(n5343), .B(n6523), .C(n5342), .D(n6518), .Q(n2321) );
  OAI222 U636 ( .A(n4851), .B(n6550), .C(n4850), .D(n6546), .Q(n2328) );
  OAI222 U637 ( .A(n4987), .B(n6541), .C(n4986), .D(n2011), .Q(n2327) );
  OAI222 U638 ( .A(n4989), .B(n6532), .C(n4988), .D(n6528), .Q(n2326) );
  OAI222 U639 ( .A(n5333), .B(n6523), .C(n5332), .D(n2015), .Q(n2325) );
  OAI222 U640 ( .A(n4609), .B(n2020), .C(n4608), .D(n2021), .Q(n2317) );
  OAI222 U641 ( .A(n4607), .B(n2022), .C(n4606), .D(n2023), .Q(n2316) );
  OAI212 U642 ( .A(n2024), .B(n5958), .C(n2329), .Q(n2315) );
  OAI222 U645 ( .A(n1162), .B(n5903), .C(n6465), .D(n5856), .Q(n2331) );
  OAI222 U646 ( .A(n4738), .B(n2032), .C(n2033), .D(n5984), .Q(n2330) );
  OAI222 U651 ( .A(n2340), .B(n6494), .C(n6316), .D(n2341), .Q(n2339) );
  OAI222 U653 ( .A(n5325), .B(n6550), .C(n5324), .D(n6546), .Q(n2345) );
  OAI222 U654 ( .A(n5183), .B(n6541), .C(n5182), .D(n6536), .Q(n2344) );
  OAI222 U655 ( .A(n5185), .B(n6532), .C(n5184), .D(n2013), .Q(n2343) );
  OAI222 U656 ( .A(n5187), .B(n6523), .C(n5186), .D(n2015), .Q(n2342) );
  OAI222 U658 ( .A(n4865), .B(n6550), .C(n4864), .D(n6545), .Q(n2349) );
  OAI222 U659 ( .A(n5023), .B(n6541), .C(n5022), .D(n2011), .Q(n2348) );
  OAI222 U660 ( .A(n5025), .B(n6532), .C(n5024), .D(n6527), .Q(n2347) );
  OAI222 U661 ( .A(n5027), .B(n6523), .C(n5026), .D(n2015), .Q(n2346) );
  OAI222 U662 ( .A(n4613), .B(n6483), .C(n4612), .D(n6485), .Q(n2338) );
  OAI222 U663 ( .A(n4611), .B(n6479), .C(n4610), .D(n6481), .Q(n2337) );
  OAI212 U664 ( .A(n6467), .B(n5957), .C(n2350), .Q(n2336) );
  OAI222 U667 ( .A(n1162), .B(n6009), .C(n2031), .D(n5888), .Q(n2352) );
  OAI222 U668 ( .A(n4762), .B(n6456), .C(n6458), .D(n5887), .Q(n2351) );
  OAI222 U673 ( .A(n2361), .B(n6494), .C(n6318), .D(n2362), .Q(n2360) );
  OAI222 U680 ( .A(n4883), .B(n6550), .C(n4882), .D(n6546), .Q(n2370) );
  OAI222 U684 ( .A(n4617), .B(n6482), .C(n4616), .D(n6484), .Q(n2359) );
  OAI212 U686 ( .A(n6466), .B(n5872), .C(n2371), .Q(n2357) );
  OAI222 U689 ( .A(n1162), .B(n5902), .C(n6465), .D(n5855), .Q(n2373) );
  OAI222 U690 ( .A(n4790), .B(n6455), .C(n6457), .D(n5886), .Q(n2372) );
  OAI222 U695 ( .A(n2382), .B(n6494), .C(n6318), .D(n2383), .Q(n2381) );
  OAI222 U702 ( .A(n4845), .B(n6550), .C(n4844), .D(n2009), .Q(n2391) );
  OAI222 U706 ( .A(n4621), .B(n2020), .C(n4620), .D(n2021), .Q(n2380) );
  OAI212 U708 ( .A(n2024), .B(n5956), .C(n2392), .Q(n2378) );
  OAI222 U711 ( .A(n1162), .B(n6008), .C(n2031), .D(n5854), .Q(n2394) );
  OAI222 U712 ( .A(n4726), .B(n2032), .C(n2033), .D(n5983), .Q(n2393) );
  OAI222 U717 ( .A(n2403), .B(n6494), .C(n6316), .D(n2404), .Q(n2402) );
  OAI222 U724 ( .A(n4859), .B(n6549), .C(n4858), .D(n6546), .Q(n2412) );
  OAI222 U728 ( .A(n4625), .B(n6483), .C(n4624), .D(n6485), .Q(n2401) );
  OAI212 U730 ( .A(n6467), .B(n5955), .C(n2413), .Q(n2399) );
  OAI222 U733 ( .A(n1162), .B(n6007), .C(n6463), .D(n5885), .Q(n2415) );
  OAI222 U734 ( .A(n4750), .B(n6456), .C(n6458), .D(n5982), .Q(n2414) );
  OAI222 U739 ( .A(n2424), .B(n6494), .C(n6318), .D(n2425), .Q(n2423) );
  OAI222 U746 ( .A(n4879), .B(n6549), .C(n4878), .D(n6545), .Q(n2433) );
  OAI222 U750 ( .A(n4629), .B(n6482), .C(n4628), .D(n6484), .Q(n2422) );
  OAI212 U752 ( .A(n6466), .B(n5871), .C(n2434), .Q(n2420) );
  OAI222 U755 ( .A(n1162), .B(n5901), .C(n6465), .D(n5853), .Q(n2436) );
  OAI222 U756 ( .A(n4782), .B(n6455), .C(n6457), .D(n5884), .Q(n2435) );
  OAI222 U761 ( .A(n2445), .B(n6494), .C(n6316), .D(n2446), .Q(n2444) );
  OAI222 U763 ( .A(n5305), .B(n6549), .C(n5304), .D(n6546), .Q(n2450) );
  OAI222 U764 ( .A(n5299), .B(n6540), .C(n5298), .D(n6536), .Q(n2449) );
  OAI222 U765 ( .A(n5301), .B(n6531), .C(n5300), .D(n6528), .Q(n2448) );
  OAI222 U766 ( .A(n5303), .B(n6522), .C(n5302), .D(n6519), .Q(n2447) );
  OAI222 U768 ( .A(n5309), .B(n6549), .C(n5308), .D(n6545), .Q(n2454) );
  OAI222 U769 ( .A(n5293), .B(n6540), .C(n5292), .D(n6536), .Q(n2453) );
  OAI222 U770 ( .A(n5295), .B(n6531), .C(n5294), .D(n6528), .Q(n2452) );
  OAI222 U771 ( .A(n5297), .B(n6522), .C(n5296), .D(n6519), .Q(n2451) );
  OAI222 U772 ( .A(n4665), .B(n2020), .C(n4664), .D(n2021), .Q(n2443) );
  OAI222 U773 ( .A(n4663), .B(n2022), .C(n4662), .D(n2023), .Q(n2442) );
  OAI212 U774 ( .A(n2024), .B(n5954), .C(n2455), .Q(n2441) );
  OAI222 U777 ( .A(n1162), .B(n6006), .C(n6460), .D(n5839), .Q(n2457) );
  OAI222 U778 ( .A(n5306), .B(n2032), .C(n2033), .D(n5981), .Q(n2456) );
  OAI222 U783 ( .A(n2466), .B(n6494), .C(n6318), .D(n2467), .Q(n2465) );
  OAI222 U790 ( .A(n4901), .B(n6549), .C(n4900), .D(n2009), .Q(n2475) );
  OAI222 U794 ( .A(n4669), .B(n6483), .C(n4668), .D(n6485), .Q(n2464) );
  OAI212 U796 ( .A(n6467), .B(n5870), .C(n2476), .Q(n2462) );
  OAI222 U799 ( .A(n1162), .B(n5900), .C(n6462), .D(n5852), .Q(n2478) );
  OAI222 U800 ( .A(n4810), .B(n6456), .C(n6458), .D(n5883), .Q(n2477) );
  OAI222 U805 ( .A(n2487), .B(n6495), .C(n6316), .D(n2488), .Q(n2486) );
  OAI222 U807 ( .A(n4891), .B(n6549), .C(n4890), .D(n6546), .Q(n2492) );
  OAI222 U808 ( .A(n5105), .B(n6540), .C(n5104), .D(n6536), .Q(n2491) );
  OAI222 U809 ( .A(n5107), .B(n6531), .C(n5106), .D(n6528), .Q(n2490) );
  OAI222 U810 ( .A(n5109), .B(n6522), .C(n5108), .D(n6519), .Q(n2489) );
  OAI222 U812 ( .A(n4847), .B(n6549), .C(n4846), .D(n2009), .Q(n2496) );
  OAI222 U813 ( .A(n4977), .B(n6540), .C(n4976), .D(n6536), .Q(n2495) );
  OAI222 U814 ( .A(n4979), .B(n6531), .C(n4978), .D(n6528), .Q(n2494) );
  OAI222 U815 ( .A(n4981), .B(n6522), .C(n4980), .D(n6519), .Q(n2493) );
  OAI222 U816 ( .A(n4673), .B(n6482), .C(n4672), .D(n6484), .Q(n2485) );
  OAI222 U817 ( .A(n4671), .B(n6478), .C(n4670), .D(n6480), .Q(n2484) );
  OAI212 U818 ( .A(n6466), .B(n5973), .C(n2497), .Q(n2483) );
  OAI222 U821 ( .A(n1162), .B(n6019), .C(n6460), .D(n5875), .Q(n2499) );
  OAI222 U822 ( .A(n4730), .B(n6455), .C(n6457), .D(n5874), .Q(n2498) );
  OAI222 U827 ( .A(n2508), .B(n6495), .C(n6316), .D(n2509), .Q(n2507) );
  OAI222 U834 ( .A(n4861), .B(n6548), .C(n4860), .D(n2009), .Q(n2517) );
  OAI222 U838 ( .A(n4677), .B(n2020), .C(n4676), .D(n2021), .Q(n2506) );
  OAI212 U840 ( .A(n2024), .B(n5869), .C(n2518), .Q(n2504) );
  OAI222 U843 ( .A(n1162), .B(n5899), .C(n6460), .D(n5851), .Q(n2520) );
  OAI222 U844 ( .A(n4754), .B(n2032), .C(n2033), .D(n5882), .Q(n2519) );
  OAI222 U849 ( .A(n2529), .B(n6495), .C(n6316), .D(n2530), .Q(n2528) );
  OAI222 U856 ( .A(n4881), .B(n6548), .C(n4880), .D(n6546), .Q(n2538) );
  OAI222 U860 ( .A(n4681), .B(n6483), .C(n4680), .D(n6485), .Q(n2527) );
  OAI212 U862 ( .A(n6467), .B(n5953), .C(n2539), .Q(n2525) );
  OAI222 U865 ( .A(n1162), .B(n6005), .C(n6464), .D(n5881), .Q(n2541) );
  OAI222 U866 ( .A(n4786), .B(n6456), .C(n6458), .D(n5980), .Q(n2540) );
  OAI222 U871 ( .A(n2550), .B(n6495), .C(n6318), .D(n2551), .Q(n2549) );
  OAI222 U878 ( .A(n4903), .B(n6548), .C(n4902), .D(n6545), .Q(n2559) );
  OAI222 U882 ( .A(n4685), .B(n6482), .C(n4684), .D(n6484), .Q(n2548) );
  OAI212 U884 ( .A(n6466), .B(n5952), .C(n2560), .Q(n2546) );
  OAI222 U887 ( .A(n1162), .B(n6004), .C(n6460), .D(n5880), .Q(n2562) );
  OAI222 U888 ( .A(n4814), .B(n6455), .C(n6457), .D(n5979), .Q(n2561) );
  OAI222 U893 ( .A(n2571), .B(n6495), .C(n6316), .D(n2572), .Q(n2570) );
  OAI222 U900 ( .A(n5347), .B(n6548), .C(n5346), .D(n6545), .Q(n2580) );
  OAI222 U904 ( .A(n4689), .B(n2020), .C(n4688), .D(n2021), .Q(n2569) );
  OAI212 U906 ( .A(n2024), .B(n5951), .C(n2581), .Q(n2567) );
  OAI222 U909 ( .A(n1162), .B(n6003), .C(n6463), .D(n5879), .Q(n2583) );
  OAI222 U910 ( .A(n4722), .B(n2032), .C(n2033), .D(n5978), .Q(n2582) );
  OAI222 U915 ( .A(n2592), .B(n6495), .C(n6318), .D(n2593), .Q(n2591) );
  OAI222 U917 ( .A(n4907), .B(n6548), .C(n4906), .D(n6545), .Q(n2597) );
  OAI222 U918 ( .A(n5151), .B(n6539), .C(n5150), .D(n6537), .Q(n2596) );
  OAI222 U919 ( .A(n5153), .B(n6530), .C(n5152), .D(n6527), .Q(n2595) );
  OAI222 U920 ( .A(n5155), .B(n6521), .C(n5154), .D(n6518), .Q(n2594) );
  OAI222 U922 ( .A(n4857), .B(n6547), .C(n4856), .D(n6545), .Q(n2601) );
  OAI222 U923 ( .A(n5001), .B(n6538), .C(n5000), .D(n6537), .Q(n2600) );
  OAI222 U925 ( .A(n5005), .B(n6520), .C(n5004), .D(n6518), .Q(n2598) );
  OAI222 U926 ( .A(n4693), .B(n6483), .C(n4692), .D(n6485), .Q(n2590) );
  OAI222 U927 ( .A(n4691), .B(n6479), .C(n4690), .D(n6481), .Q(n2589) );
  OAI212 U928 ( .A(n6467), .B(n5972), .C(n2602), .Q(n2588) );
  OAI222 U931 ( .A(n1162), .B(n6018), .C(n6460), .D(n5897), .Q(n2604) );
  OAI222 U932 ( .A(n4746), .B(n6456), .C(n6458), .D(n5998), .Q(n2603) );
  OAI222 U937 ( .A(n2613), .B(n6495), .C(n6316), .D(n2614), .Q(n2612) );
  OAI222 U944 ( .A(n4875), .B(n6547), .C(n4874), .D(n6545), .Q(n2622) );
  OAI222 U948 ( .A(n4697), .B(n6482), .C(n4696), .D(n6484), .Q(n2611) );
  OAI212 U950 ( .A(n6466), .B(n5950), .C(n2623), .Q(n2609) );
  OAI222 U953 ( .A(n1162), .B(n6002), .C(n6462), .D(n5878), .Q(n2625) );
  OAI222 U954 ( .A(n4778), .B(n6455), .C(n6457), .D(n5977), .Q(n2624) );
  OAI222 U959 ( .A(n2634), .B(n6495), .C(n6316), .D(n2635), .Q(n2633) );
  OAI222 U966 ( .A(n4893), .B(n6547), .C(n4892), .D(n6545), .Q(n2643) );
  OAI222 U970 ( .A(n4701), .B(n2020), .C(n4700), .D(n2021), .Q(n2632) );
  OAI212 U972 ( .A(n2024), .B(n5949), .C(n2644), .Q(n2630) );
  OAI222 U975 ( .A(n1162), .B(n6001), .C(n6460), .D(n5877), .Q(n2646) );
  OAI222 U976 ( .A(n4802), .B(n2032), .C(n2033), .D(n5976), .Q(n2645) );
  OAI222 U981 ( .A(n2655), .B(n6495), .C(n6316), .D(n2656), .Q(n2654) );
  OAI222 U988 ( .A(n4855), .B(n6547), .C(n4854), .D(n6545), .Q(n2664) );
  OAI222 U992 ( .A(n4705), .B(n6483), .C(n4704), .D(n6485), .Q(n2653) );
  OAI212 U994 ( .A(n6467), .B(n5948), .C(n2665), .Q(n2651) );
  OAI222 U997 ( .A(n1162), .B(n6000), .C(n6462), .D(n5876), .Q(n2667) );
  OAI222 U998 ( .A(n4742), .B(n6456), .C(n6458), .D(n5975), .Q(n2666) );
  OAI222 U1003 ( .A(n2676), .B(n6492), .C(n6316), .D(n2677), .Q(n2675) );
  OAI222 U1005 ( .A(n5331), .B(n6547), .C(n5330), .D(n6545), .Q(n2681) );
  OAI222 U1006 ( .A(n5287), .B(n6538), .C(n5286), .D(n6537), .Q(n2680) );
  OAI222 U1007 ( .A(n5289), .B(n6529), .C(n5288), .D(n6527), .Q(n2679) );
  OAI222 U1008 ( .A(n5291), .B(n6520), .C(n5290), .D(n6518), .Q(n2678) );
  OAI222 U1010 ( .A(n4837), .B(n6547), .C(n4836), .D(n6545), .Q(n2685) );
  OAI222 U1013 ( .A(n4949), .B(n6538), .C(n4948), .D(n6536), .Q(n2684) );
  OAI222 U1020 ( .A(n5315), .B(n6520), .C(n5314), .D(n6518), .Q(n2682) );
  OAI222 U1024 ( .A(n4709), .B(n6482), .C(n4708), .D(n6484), .Q(n2674) );
  OAI222 U1027 ( .A(n4707), .B(n6478), .C(n4706), .D(n6480), .Q(n2673) );
  OAI212 U1030 ( .A(n6466), .B(n5947), .C(n2695), .Q(n2672) );
  OAI222 U1036 ( .A(n1162), .B(n5898), .C(n5692), .D(n6465), .Q(n2699) );
  OAI222 U1040 ( .A(n4830), .B(n6455), .C(n6457), .D(n5974), .Q(n2698) );
  OAI222 U1065 ( .A(n2714), .B(n6499), .C(n6320), .D(n2715), .Q(n2713) );
  OAI222 U1067 ( .A(n5319), .B(n6590), .C(n5318), .D(n1926), .Q(n2719) );
  OAI222 U1068 ( .A(n5201), .B(n6580), .C(n5200), .D(n1928), .Q(n2718) );
  OAI222 U1069 ( .A(n5203), .B(n6571), .C(n5202), .D(n6564), .Q(n2717) );
  OAI222 U1070 ( .A(n5205), .B(n6562), .C(n5204), .D(n1932), .Q(n2716) );
  OAI222 U1072 ( .A(n4873), .B(n6590), .C(n4872), .D(n6582), .Q(n2723) );
  OAI222 U1073 ( .A(n5047), .B(n6580), .C(n5046), .D(n1928), .Q(n2722) );
  OAI222 U1074 ( .A(n5049), .B(n6571), .C(n5048), .D(n6564), .Q(n2721) );
  OAI222 U1075 ( .A(n5341), .B(n6562), .C(n5340), .D(n1932), .Q(n2720) );
  OAI222 U1076 ( .A(n4633), .B(n6418), .C(n4632), .D(n6420), .Q(n2712) );
  OAI222 U1077 ( .A(n4631), .B(n6414), .C(n4630), .D(n6416), .Q(n2711) );
  OAI212 U1078 ( .A(n1941), .B(n5971), .C(n2724), .Q(n2710) );
  OAI222 U1081 ( .A(n1170), .B(n6017), .C(n6400), .D(n5857), .Q(n2726) );
  OAI222 U1082 ( .A(n4774), .B(n6392), .C(n1950), .D(n5997), .Q(n2725) );
  OAI222 U1087 ( .A(n2735), .B(n6499), .C(n6320), .D(n2736), .Q(n2734) );
  OAI222 U1089 ( .A(n4939), .B(n6590), .C(n4938), .D(n6581), .Q(n2740) );
  OAI222 U1090 ( .A(n5253), .B(n6580), .C(n5252), .D(n1928), .Q(n2739) );
  OAI222 U1091 ( .A(n5255), .B(n6571), .C(n5254), .D(n6564), .Q(n2738) );
  OAI222 U1092 ( .A(n5257), .B(n6562), .C(n5256), .D(n1932), .Q(n2737) );
  OAI222 U1094 ( .A(n4897), .B(n6590), .C(n4896), .D(n6581), .Q(n2744) );
  OAI222 U1095 ( .A(n5123), .B(n6580), .C(n5122), .D(n1928), .Q(n2743) );
  OAI222 U1096 ( .A(n5125), .B(n6571), .C(n5124), .D(n6564), .Q(n2742) );
  OAI222 U1098 ( .A(n4637), .B(n1937), .C(n4636), .D(n1938), .Q(n2733) );
  OAI222 U1099 ( .A(n4635), .B(n1939), .C(n4634), .D(n1940), .Q(n2732) );
  OAI212 U1100 ( .A(n6403), .B(n5970), .C(n2745), .Q(n2731) );
  OAI222 U1103 ( .A(n1170), .B(n6016), .C(n1948), .D(n5896), .Q(n2747) );
  OAI222 U1104 ( .A(n4806), .B(n1949), .C(n6396), .D(n5996), .Q(n2746) );
  OAI222 U1109 ( .A(n2756), .B(n6499), .C(n6319), .D(n2757), .Q(n2755) );
  OAI222 U1111 ( .A(n4947), .B(n6590), .C(n4946), .D(n1926), .Q(n2761) );
  OAI222 U1112 ( .A(n5275), .B(n6580), .C(n5274), .D(n1928), .Q(n2760) );
  OAI222 U1113 ( .A(n5277), .B(n6571), .C(n5276), .D(n6564), .Q(n2759) );
  OAI222 U1114 ( .A(n5279), .B(n6562), .C(n5278), .D(n1932), .Q(n2758) );
  OAI222 U1116 ( .A(n4917), .B(n6590), .C(n4916), .D(n1926), .Q(n2765) );
  OAI222 U1117 ( .A(n5177), .B(n6580), .C(n5176), .D(n1928), .Q(n2764) );
  OAI222 U1118 ( .A(n5179), .B(n6571), .C(n5178), .D(n6564), .Q(n2763) );
  OAI222 U1119 ( .A(n5181), .B(n6562), .C(n5180), .D(n1932), .Q(n2762) );
  OAI222 U1120 ( .A(n4641), .B(n6419), .C(n4640), .D(n6421), .Q(n2754) );
  OAI222 U1121 ( .A(n4639), .B(n6415), .C(n4638), .D(n6417), .Q(n2753) );
  OAI212 U1122 ( .A(n6402), .B(n5969), .C(n2766), .Q(n2752) );
  OAI222 U1125 ( .A(n1170), .B(n6015), .C(n6401), .D(n5895), .Q(n2768) );
  OAI222 U1126 ( .A(n4822), .B(n6393), .C(n6396), .D(n5995), .Q(n2767) );
  OAI222 U1131 ( .A(n2777), .B(n6499), .C(n6319), .D(n2778), .Q(n2776) );
  OAI222 U1133 ( .A(n4919), .B(n6590), .C(n4918), .D(n1926), .Q(n2782) );
  OAI222 U1134 ( .A(n5189), .B(n6580), .C(n5188), .D(n6572), .Q(n2781) );
  OAI222 U1135 ( .A(n5191), .B(n6571), .C(n5190), .D(n6564), .Q(n2780) );
  OAI222 U1136 ( .A(n5193), .B(n6562), .C(n5192), .D(n1932), .Q(n2779) );
  OAI222 U1138 ( .A(n4867), .B(n6590), .C(n4866), .D(n1926), .Q(n2786) );
  OAI222 U1139 ( .A(n5029), .B(n6580), .C(n5028), .D(n1928), .Q(n2785) );
  OAI222 U1140 ( .A(n5031), .B(n6571), .C(n5030), .D(n6564), .Q(n2784) );
  OAI222 U1141 ( .A(n5033), .B(n6562), .C(n5032), .D(n1932), .Q(n2783) );
  OAI222 U1142 ( .A(n4645), .B(n6418), .C(n4644), .D(n6420), .Q(n2775) );
  OAI222 U1143 ( .A(n4643), .B(n6414), .C(n4642), .D(n6416), .Q(n2774) );
  OAI212 U1144 ( .A(n1941), .B(n5968), .C(n2787), .Q(n2773) );
  OAI222 U1147 ( .A(n1170), .B(n6014), .C(n6400), .D(n5894), .Q(n2789) );
  OAI222 U1148 ( .A(n4766), .B(n6392), .C(n6397), .D(n5994), .Q(n2788) );
  OAI222 U1153 ( .A(n2798), .B(n6499), .C(n6319), .D(n2799), .Q(n2797) );
  OAI222 U1155 ( .A(n4933), .B(n6589), .C(n4932), .D(n1926), .Q(n2803) );
  OAI222 U1156 ( .A(n5235), .B(n6579), .C(n5234), .D(n6573), .Q(n2802) );
  OAI222 U1157 ( .A(n5237), .B(n6570), .C(n5236), .D(n6564), .Q(n2801) );
  OAI222 U1158 ( .A(n5239), .B(n6561), .C(n5238), .D(n6554), .Q(n2800) );
  OAI222 U1160 ( .A(n4887), .B(n6589), .C(n4886), .D(n1926), .Q(n2807) );
  OAI222 U1161 ( .A(n5087), .B(n6579), .C(n5086), .D(n6573), .Q(n2806) );
  OAI222 U1162 ( .A(n5089), .B(n6570), .C(n5088), .D(n6564), .Q(n2805) );
  OAI222 U1163 ( .A(n5091), .B(n6561), .C(n5090), .D(n1932), .Q(n2804) );
  OAI222 U1164 ( .A(n4649), .B(n1937), .C(n4648), .D(n1938), .Q(n2796) );
  OAI222 U1165 ( .A(n4647), .B(n1939), .C(n4646), .D(n1940), .Q(n2795) );
  OAI212 U1166 ( .A(n6403), .B(n5967), .C(n2808), .Q(n2794) );
  OAI222 U1169 ( .A(n1170), .B(n6013), .C(n1948), .D(n5893), .Q(n2810) );
  OAI222 U1170 ( .A(n4794), .B(n1949), .C(n6398), .D(n5993), .Q(n2809) );
  OAI222 U1175 ( .A(n2819), .B(n6499), .C(n6319), .D(n2820), .Q(n2818) );
  OAI222 U1177 ( .A(n4945), .B(n6589), .C(n4944), .D(n1926), .Q(n2824) );
  OAI222 U1178 ( .A(n5271), .B(n6579), .C(n5270), .D(n1928), .Q(n2823) );
  OAI222 U1179 ( .A(n5273), .B(n6570), .C(n5272), .D(n6564), .Q(n2822) );
  OAI222 U1180 ( .A(n5345), .B(n6561), .C(n5344), .D(n1932), .Q(n2821) );
  OAI222 U1182 ( .A(n4909), .B(n6589), .C(n4908), .D(n1926), .Q(n2828) );
  OAI222 U1183 ( .A(n5157), .B(n6579), .C(n5156), .D(n1928), .Q(n2827) );
  OAI222 U1184 ( .A(n5159), .B(n6570), .C(n5158), .D(n6563), .Q(n2826) );
  OAI222 U1185 ( .A(n5327), .B(n6561), .C(n5326), .D(n1932), .Q(n2825) );
  OAI222 U1186 ( .A(n4653), .B(n6419), .C(n4652), .D(n6421), .Q(n2817) );
  OAI222 U1187 ( .A(n4651), .B(n6415), .C(n4650), .D(n6417), .Q(n2816) );
  OAI212 U1188 ( .A(n6402), .B(n5966), .C(n2829), .Q(n2815) );
  OAI222 U1191 ( .A(n1170), .B(n6012), .C(n6401), .D(n5892), .Q(n2831) );
  OAI222 U1192 ( .A(n4818), .B(n6393), .C(n6398), .D(n5992), .Q(n2830) );
  OAI222 U1197 ( .A(n2840), .B(n6499), .C(n6319), .D(n2841), .Q(n2839) );
  OAI222 U1199 ( .A(n5321), .B(n6589), .C(n5320), .D(n1926), .Q(n2845) );
  OAI222 U1200 ( .A(n5281), .B(n6579), .C(n5280), .D(n1928), .Q(n2844) );
  OAI222 U1201 ( .A(n5283), .B(n6570), .C(n5282), .D(n6564), .Q(n2843) );
  OAI222 U1202 ( .A(n5285), .B(n6561), .C(n5284), .D(n1932), .Q(n2842) );
  OAI222 U1204 ( .A(n4925), .B(n6589), .C(n4924), .D(n1926), .Q(n2849) );
  OAI222 U1205 ( .A(n5213), .B(n6579), .C(n5212), .D(n1928), .Q(n2848) );
  OAI222 U1206 ( .A(n5215), .B(n6570), .C(n5214), .D(n6563), .Q(n2847) );
  OAI222 U1207 ( .A(n5317), .B(n6561), .C(n5316), .D(n1932), .Q(n2846) );
  OAI222 U1208 ( .A(n4657), .B(n6418), .C(n4656), .D(n6420), .Q(n2838) );
  OAI222 U1209 ( .A(n4655), .B(n6414), .C(n4654), .D(n6416), .Q(n2837) );
  OAI212 U1210 ( .A(n1941), .B(n5965), .C(n2850), .Q(n2836) );
  OAI222 U1213 ( .A(n1170), .B(n6011), .C(n6400), .D(n5891), .Q(n2852) );
  OAI222 U1214 ( .A(n4826), .B(n6392), .C(n6399), .D(n5991), .Q(n2851) );
  OAI222 U1219 ( .A(n2861), .B(n6499), .C(n6319), .D(n2862), .Q(n2860) );
  OAI222 U1224 ( .A(n5245), .B(n6561), .C(n5244), .D(n1932), .Q(n2863) );
  OAI222 U1226 ( .A(n4889), .B(n6589), .C(n4888), .D(n1926), .Q(n2870) );
  OAI222 U1230 ( .A(n4585), .B(n1937), .C(n4584), .D(n1938), .Q(n2859) );
  OAI212 U1232 ( .A(n6403), .B(n5873), .C(n2871), .Q(n2857) );
  OAI222 U1236 ( .A(n4798), .B(n1949), .C(n1950), .D(n5890), .Q(n2872) );
  OAI222 U1241 ( .A(n2882), .B(n6500), .C(n6319), .D(n2883), .Q(n2881) );
  OAI222 U1244 ( .A(n4991), .B(n6579), .C(n4990), .D(n6573), .Q(n2886) );
  OAI222 U1245 ( .A(n4993), .B(n6570), .C(n4992), .D(n1930), .Q(n2885) );
  OAI222 U1246 ( .A(n4995), .B(n6561), .C(n4994), .D(n6555), .Q(n2884) );
  OAI222 U1248 ( .A(n4839), .B(n6588), .C(n4838), .D(n1926), .Q(n2891) );
  OAI222 U1250 ( .A(n4955), .B(n6569), .C(n4954), .D(n6564), .Q(n2889) );
  OAI222 U1251 ( .A(n4957), .B(n6560), .C(n4956), .D(n6554), .Q(n2888) );
  OAI222 U1252 ( .A(n4589), .B(n6419), .C(n4588), .D(n6421), .Q(n2880) );
  OAI212 U1254 ( .A(n6402), .B(n5964), .C(n2892), .Q(n2878) );
  OAI222 U1257 ( .A(n1170), .B(n6062), .C(n6401), .D(n5904), .Q(n2894) );
  OAI222 U1258 ( .A(n4710), .B(n6393), .C(n1950), .D(n5990), .Q(n2893) );
  OAI222 U1263 ( .A(n2903), .B(n6499), .C(n6319), .D(n2904), .Q(n2902) );
  OAI222 U1267 ( .A(n5197), .B(n6569), .C(n5196), .D(n1930), .Q(n2906) );
  OAI222 U1268 ( .A(n5199), .B(n6560), .C(n5198), .D(n1932), .Q(n2905) );
  OAI222 U1270 ( .A(n4869), .B(n6588), .C(n4868), .D(n1926), .Q(n2912) );
  OAI222 U1274 ( .A(n4661), .B(n6418), .C(n4660), .D(n6420), .Q(n2901) );
  OAI212 U1276 ( .A(n1941), .B(n5963), .C(n2913), .Q(n2899) );
  OAI222 U1280 ( .A(n4770), .B(n6392), .C(n1950), .D(n5989), .Q(n2914) );
  OAI222 U1285 ( .A(n2924), .B(n6499), .C(n6320), .D(n2925), .Q(n2923) );
  OAI222 U1289 ( .A(n5043), .B(n6569), .C(n5042), .D(n6564), .Q(n2927) );
  OAI222 U1290 ( .A(n5045), .B(n6560), .C(n5044), .D(n1932), .Q(n2926) );
  OAI222 U1292 ( .A(n4841), .B(n6588), .C(n4840), .D(n1926), .Q(n2933) );
  OAI222 U1296 ( .A(n4593), .B(n1937), .C(n4592), .D(n1938), .Q(n2922) );
  OAI212 U1298 ( .A(n6403), .B(n5962), .C(n2934), .Q(n2920) );
  OAI222 U1302 ( .A(n4714), .B(n1949), .C(n6399), .D(n5988), .Q(n2935) );
  OAI222 U1307 ( .A(n2945), .B(n6500), .C(n6319), .D(n2946), .Q(n2944) );
  OAI222 U1311 ( .A(n5119), .B(n6569), .C(n5118), .D(n6564), .Q(n2948) );
  OAI222 U1312 ( .A(n5121), .B(n6560), .C(n5120), .D(n1932), .Q(n2947) );
  OAI222 U1314 ( .A(n4849), .B(n6588), .C(n4848), .D(n6583), .Q(n2954) );
  OAI222 U1318 ( .A(n4597), .B(n6419), .C(n4596), .D(n6421), .Q(n2943) );
  OAI212 U1320 ( .A(n6402), .B(n5961), .C(n2955), .Q(n2941) );
  OAI222 U1324 ( .A(n4734), .B(n6393), .C(n6397), .D(n5987), .Q(n2956) );
  OAI222 U1329 ( .A(n2966), .B(n6500), .C(n6319), .D(n2967), .Q(n2965) );
  OAI222 U1331 ( .A(n4915), .B(n6588), .C(n4914), .D(n6583), .Q(n2971) );
  OAI222 U1332 ( .A(n5173), .B(n6578), .C(n5172), .D(n6573), .Q(n2970) );
  OAI222 U1333 ( .A(n5175), .B(n6569), .C(n5174), .D(n6563), .Q(n2969) );
  OAI222 U1334 ( .A(n5335), .B(n6560), .C(n5334), .D(n6555), .Q(n2968) );
  OAI222 U1336 ( .A(n4863), .B(n6588), .C(n4862), .D(n6583), .Q(n2975) );
  OAI222 U1337 ( .A(n5017), .B(n6578), .C(n5016), .D(n6573), .Q(n2974) );
  OAI222 U1338 ( .A(n5019), .B(n6569), .C(n5018), .D(n1930), .Q(n2973) );
  OAI222 U1339 ( .A(n5021), .B(n6560), .C(n5020), .D(n6555), .Q(n2972) );
  OAI222 U1340 ( .A(n4601), .B(n6418), .C(n4600), .D(n6420), .Q(n2964) );
  OAI222 U1341 ( .A(n4599), .B(n6414), .C(n4598), .D(n6416), .Q(n2963) );
  OAI212 U1342 ( .A(n1941), .B(n5960), .C(n2976), .Q(n2962) );
  OAI222 U1345 ( .A(n1170), .B(n6010), .C(n6400), .D(n5889), .Q(n2978) );
  OAI222 U1346 ( .A(n4758), .B(n6392), .C(n6396), .D(n5986), .Q(n2977) );
  OAI222 U1351 ( .A(n2987), .B(n6500), .C(n6319), .D(n2988), .Q(n2986) );
  OAI222 U1353 ( .A(n4877), .B(n6587), .C(n4876), .D(n6583), .Q(n2992) );
  OAI222 U1354 ( .A(n5057), .B(n6577), .C(n5056), .D(n6573), .Q(n2991) );
  OAI222 U1355 ( .A(n5059), .B(n6568), .C(n5058), .D(n1930), .Q(n2990) );
  OAI222 U1356 ( .A(n5061), .B(n6559), .C(n5060), .D(n6555), .Q(n2989) );
  OAI222 U1359 ( .A(n4965), .B(n6577), .C(n4964), .D(n6573), .Q(n2995) );
  OAI222 U1360 ( .A(n4967), .B(n6568), .C(n4966), .D(n1930), .Q(n2994) );
  OAI222 U1361 ( .A(n5339), .B(n6559), .C(n5338), .D(n6555), .Q(n2993) );
  OAI222 U1362 ( .A(n4605), .B(n1937), .C(n4604), .D(n1938), .Q(n2985) );
  OAI212 U1364 ( .A(n6403), .B(n5959), .C(n2997), .Q(n2983) );
  OAI222 U1368 ( .A(n4718), .B(n1949), .C(n1950), .D(n5985), .Q(n2998) );
  OAI222 U1373 ( .A(n3008), .B(n6500), .C(n6319), .D(n3009), .Q(n3007) );
  OAI222 U1375 ( .A(n4899), .B(n6587), .C(n4898), .D(n6583), .Q(n3013) );
  OAI222 U1376 ( .A(n5129), .B(n6577), .C(n5128), .D(n6573), .Q(n3012) );
  OAI222 U1377 ( .A(n5131), .B(n6568), .C(n5130), .D(n1930), .Q(n3011) );
  OAI222 U1378 ( .A(n5343), .B(n6559), .C(n5342), .D(n6555), .Q(n3010) );
  OAI222 U1380 ( .A(n4851), .B(n6587), .C(n4850), .D(n6583), .Q(n3017) );
  OAI222 U1381 ( .A(n4987), .B(n6577), .C(n4986), .D(n6573), .Q(n3016) );
  OAI222 U1382 ( .A(n4989), .B(n6568), .C(n4988), .D(n1930), .Q(n3015) );
  OAI222 U1383 ( .A(n5333), .B(n6559), .C(n5332), .D(n6555), .Q(n3014) );
  OAI222 U1384 ( .A(n4609), .B(n6419), .C(n4608), .D(n6421), .Q(n3006) );
  OAI222 U1385 ( .A(n4607), .B(n6415), .C(n4606), .D(n6417), .Q(n3005) );
  OAI212 U1386 ( .A(n6402), .B(n5958), .C(n3018), .Q(n3004) );
  OAI222 U1389 ( .A(n1170), .B(n5903), .C(n6401), .D(n5856), .Q(n3020) );
  OAI222 U1390 ( .A(n4738), .B(n6393), .C(n1950), .D(n5984), .Q(n3019) );
  OAI222 U1395 ( .A(n3029), .B(n6500), .C(n6319), .D(n3030), .Q(n3028) );
  OAI222 U1397 ( .A(n5325), .B(n6587), .C(n5324), .D(n6583), .Q(n3034) );
  OAI222 U1398 ( .A(n5183), .B(n6577), .C(n5182), .D(n6573), .Q(n3033) );
  OAI222 U1399 ( .A(n5185), .B(n6568), .C(n5184), .D(n1930), .Q(n3032) );
  OAI222 U1400 ( .A(n5187), .B(n6559), .C(n5186), .D(n6555), .Q(n3031) );
  OAI222 U1402 ( .A(n4865), .B(n6587), .C(n4864), .D(n6583), .Q(n3038) );
  OAI222 U1403 ( .A(n5023), .B(n6577), .C(n5022), .D(n6573), .Q(n3037) );
  OAI222 U1404 ( .A(n5025), .B(n6568), .C(n5024), .D(n1930), .Q(n3036) );
  OAI222 U1405 ( .A(n5027), .B(n6559), .C(n5026), .D(n6555), .Q(n3035) );
  OAI222 U1406 ( .A(n4613), .B(n6418), .C(n4612), .D(n6420), .Q(n3027) );
  OAI222 U1407 ( .A(n4611), .B(n6414), .C(n4610), .D(n6416), .Q(n3026) );
  OAI212 U1408 ( .A(n1941), .B(n5957), .C(n3039), .Q(n3025) );
  OAI222 U1411 ( .A(n1170), .B(n6009), .C(n6400), .D(n5888), .Q(n3041) );
  OAI222 U1412 ( .A(n4762), .B(n6392), .C(n6399), .D(n5887), .Q(n3040) );
  OAI222 U1417 ( .A(n3050), .B(n6500), .C(n6319), .D(n3051), .Q(n3049) );
  OAI222 U1419 ( .A(n4931), .B(n6587), .C(n4930), .D(n6583), .Q(n3055) );
  OAI222 U1420 ( .A(n5229), .B(n6577), .C(n5228), .D(n6573), .Q(n3054) );
  OAI222 U1421 ( .A(n5231), .B(n6568), .C(n5230), .D(n1930), .Q(n3053) );
  OAI222 U1422 ( .A(n5233), .B(n6559), .C(n5232), .D(n6555), .Q(n3052) );
  OAI222 U1424 ( .A(n4883), .B(n6587), .C(n4882), .D(n6583), .Q(n3059) );
  OAI222 U1425 ( .A(n5075), .B(n6577), .C(n5074), .D(n6573), .Q(n3058) );
  OAI222 U1426 ( .A(n5077), .B(n6568), .C(n5076), .D(n1930), .Q(n3057) );
  OAI222 U1427 ( .A(n5079), .B(n6559), .C(n5078), .D(n6555), .Q(n3056) );
  OAI222 U1428 ( .A(n4617), .B(n1937), .C(n4616), .D(n1938), .Q(n3048) );
  OAI222 U1429 ( .A(n4615), .B(n1939), .C(n4614), .D(n1940), .Q(n3047) );
  OAI212 U1430 ( .A(n6403), .B(n5872), .C(n3060), .Q(n3046) );
  OAI222 U1433 ( .A(n1170), .B(n5902), .C(n1948), .D(n5855), .Q(n3062) );
  OAI222 U1434 ( .A(n4790), .B(n1949), .C(n6399), .D(n5886), .Q(n3061) );
  OAI222 U1439 ( .A(n3071), .B(n6500), .C(n6319), .D(n3072), .Q(n3070) );
  OAI222 U1441 ( .A(n5329), .B(n6587), .C(n5328), .D(n6583), .Q(n3076) );
  OAI222 U1442 ( .A(n5093), .B(n6577), .C(n5092), .D(n6573), .Q(n3075) );
  OAI222 U1443 ( .A(n5095), .B(n6568), .C(n5094), .D(n6563), .Q(n3074) );
  OAI222 U1444 ( .A(n5097), .B(n6559), .C(n5096), .D(n6555), .Q(n3073) );
  OAI222 U1446 ( .A(n4845), .B(n6586), .C(n4844), .D(n6583), .Q(n3080) );
  OAI222 U1447 ( .A(n4973), .B(n6576), .C(n4972), .D(n6573), .Q(n3079) );
  OAI222 U1448 ( .A(n4975), .B(n6567), .C(n4974), .D(n1930), .Q(n3078) );
  OAI222 U1449 ( .A(n5337), .B(n6558), .C(n5336), .D(n6555), .Q(n3077) );
  OAI222 U1450 ( .A(n4621), .B(n6419), .C(n4620), .D(n6421), .Q(n3069) );
  OAI222 U1451 ( .A(n4619), .B(n6415), .C(n4618), .D(n6417), .Q(n3068) );
  OAI212 U1452 ( .A(n6402), .B(n5956), .C(n3081), .Q(n3067) );
  OAI222 U1455 ( .A(n1170), .B(n6008), .C(n6401), .D(n5854), .Q(n3083) );
  OAI222 U1456 ( .A(n4726), .B(n6393), .C(n1950), .D(n5983), .Q(n3082) );
  OAI222 U1461 ( .A(n3092), .B(n6500), .C(n6319), .D(n3093), .Q(n3091) );
  OAI222 U1463 ( .A(n4911), .B(n6586), .C(n4910), .D(n6582), .Q(n3097) );
  OAI222 U1464 ( .A(n5161), .B(n6576), .C(n5160), .D(n6572), .Q(n3096) );
  OAI222 U1465 ( .A(n5163), .B(n6567), .C(n5162), .D(n6563), .Q(n3095) );
  OAI222 U1466 ( .A(n5165), .B(n6558), .C(n5164), .D(n6554), .Q(n3094) );
  OAI222 U1468 ( .A(n4859), .B(n6586), .C(n4858), .D(n6582), .Q(n3101) );
  OAI222 U1469 ( .A(n5007), .B(n6576), .C(n5006), .D(n1928), .Q(n3100) );
  OAI222 U1470 ( .A(n5009), .B(n6567), .C(n5008), .D(n6563), .Q(n3099) );
  OAI222 U1471 ( .A(n5323), .B(n6558), .C(n5322), .D(n6554), .Q(n3098) );
  OAI222 U1472 ( .A(n4625), .B(n6418), .C(n4624), .D(n6420), .Q(n3090) );
  OAI222 U1473 ( .A(n4623), .B(n6414), .C(n4622), .D(n6416), .Q(n3089) );
  OAI212 U1474 ( .A(n1941), .B(n5955), .C(n3102), .Q(n3088) );
  OAI222 U1477 ( .A(n1170), .B(n6007), .C(n6400), .D(n5885), .Q(n3104) );
  OAI222 U1478 ( .A(n4750), .B(n6392), .C(n1950), .D(n5982), .Q(n3103) );
  OAI222 U1483 ( .A(n3113), .B(n6500), .C(n6320), .D(n3114), .Q(n3112) );
  OAI222 U1485 ( .A(n4927), .B(n6586), .C(n4926), .D(n6582), .Q(n3118) );
  OAI222 U1486 ( .A(n5217), .B(n6576), .C(n5216), .D(n6572), .Q(n3117) );
  OAI222 U1487 ( .A(n5219), .B(n6567), .C(n5218), .D(n6563), .Q(n3116) );
  OAI222 U1488 ( .A(n5221), .B(n6558), .C(n5220), .D(n6554), .Q(n3115) );
  OAI222 U1490 ( .A(n4879), .B(n6586), .C(n4878), .D(n6582), .Q(n3122) );
  OAI222 U1491 ( .A(n5063), .B(n6576), .C(n5062), .D(n6572), .Q(n3121) );
  OAI222 U1492 ( .A(n5065), .B(n6567), .C(n5064), .D(n6563), .Q(n3120) );
  OAI222 U1493 ( .A(n5067), .B(n6558), .C(n5066), .D(n6554), .Q(n3119) );
  OAI222 U1494 ( .A(n4629), .B(n1937), .C(n4628), .D(n1938), .Q(n3111) );
  OAI222 U1495 ( .A(n4627), .B(n1939), .C(n4626), .D(n1940), .Q(n3110) );
  OAI212 U1496 ( .A(n6403), .B(n5871), .C(n3123), .Q(n3109) );
  OAI222 U1499 ( .A(n1170), .B(n5901), .C(n1948), .D(n5853), .Q(n3125) );
  OAI222 U1500 ( .A(n4782), .B(n1949), .C(n6398), .D(n5884), .Q(n3124) );
  OAI222 U1505 ( .A(n3134), .B(n6500), .C(n6319), .D(n3135), .Q(n3133) );
  OAI222 U1512 ( .A(n5309), .B(n6586), .C(n5308), .D(n6582), .Q(n3143) );
  OAI222 U1516 ( .A(n4665), .B(n6419), .C(n4664), .D(n6421), .Q(n3132) );
  OAI212 U1518 ( .A(n6402), .B(n5954), .C(n3144), .Q(n3130) );
  OAI222 U1521 ( .A(n1170), .B(n6006), .C(n6401), .D(n5839), .Q(n3146) );
  OAI222 U1522 ( .A(n5306), .B(n6393), .C(n6397), .D(n5981), .Q(n3145) );
  OAI222 U1527 ( .A(n3155), .B(n6501), .C(n6320), .D(n3156), .Q(n3154) );
  OAI222 U1529 ( .A(n4941), .B(n6586), .C(n4940), .D(n6582), .Q(n3160) );
  OAI222 U1530 ( .A(n5259), .B(n6576), .C(n5258), .D(n6573), .Q(n3159) );
  OAI222 U1531 ( .A(n5261), .B(n6567), .C(n5260), .D(n6563), .Q(n3158) );
  OAI222 U1532 ( .A(n5263), .B(n6558), .C(n5262), .D(n6554), .Q(n3157) );
  OAI222 U1534 ( .A(n4901), .B(n6586), .C(n4900), .D(n6582), .Q(n3164) );
  OAI222 U1535 ( .A(n5133), .B(n6576), .C(n5132), .D(n6573), .Q(n3163) );
  OAI222 U1536 ( .A(n5135), .B(n6567), .C(n5134), .D(n6563), .Q(n3162) );
  OAI222 U1537 ( .A(n5137), .B(n6558), .C(n5136), .D(n6554), .Q(n3161) );
  OAI222 U1538 ( .A(n4669), .B(n6418), .C(n4668), .D(n6420), .Q(n3153) );
  OAI222 U1539 ( .A(n4667), .B(n6414), .C(n4666), .D(n6416), .Q(n3152) );
  OAI212 U1540 ( .A(n1941), .B(n5870), .C(n3165), .Q(n3151) );
  OAI222 U1543 ( .A(n1170), .B(n5900), .C(n6400), .D(n5852), .Q(n3167) );
  OAI222 U1544 ( .A(n4810), .B(n6392), .C(n6397), .D(n5883), .Q(n3166) );
  OAI222 U1549 ( .A(n3176), .B(n6501), .C(n6320), .D(n3177), .Q(n3175) );
  OAI222 U1556 ( .A(n4847), .B(n6585), .C(n4846), .D(n6582), .Q(n3185) );
  OAI222 U1560 ( .A(n4673), .B(n1937), .C(n4672), .D(n1938), .Q(n3174) );
  OAI212 U1562 ( .A(n5973), .B(n6403), .C(n3186), .Q(n3172) );
  OAI222 U1565 ( .A(n6019), .B(n1170), .C(n5875), .D(n6401), .Q(n3188) );
  OAI222 U1566 ( .A(n4730), .B(n1949), .C(n5874), .D(n6399), .Q(n3187) );
  OAI222 U1571 ( .A(n3197), .B(n6501), .C(n6320), .D(n3198), .Q(n3196) );
  OAI222 U1573 ( .A(n4913), .B(n6585), .C(n4912), .D(n6582), .Q(n3202) );
  OAI222 U1574 ( .A(n5167), .B(n6575), .C(n5166), .D(n6573), .Q(n3201) );
  OAI222 U1575 ( .A(n5169), .B(n6566), .C(n5168), .D(n6563), .Q(n3200) );
  OAI222 U1576 ( .A(n5171), .B(n6557), .C(n5170), .D(n6554), .Q(n3199) );
  OAI222 U1578 ( .A(n4861), .B(n6585), .C(n4860), .D(n6582), .Q(n3206) );
  OAI222 U1579 ( .A(n5011), .B(n6575), .C(n5010), .D(n6572), .Q(n3205) );
  OAI222 U1580 ( .A(n5013), .B(n6566), .C(n5012), .D(n6563), .Q(n3204) );
  OAI222 U1581 ( .A(n5015), .B(n6557), .C(n5014), .D(n6554), .Q(n3203) );
  OAI222 U1582 ( .A(n4677), .B(n6419), .C(n4676), .D(n6421), .Q(n3195) );
  OAI222 U1583 ( .A(n4675), .B(n6415), .C(n4674), .D(n6417), .Q(n3194) );
  OAI212 U1584 ( .A(n6403), .B(n5869), .C(n3207), .Q(n3193) );
  OAI222 U1587 ( .A(n1170), .B(n5899), .C(n1948), .D(n5851), .Q(n3209) );
  OAI222 U1588 ( .A(n4754), .B(n6393), .C(n6396), .D(n5882), .Q(n3208) );
  OAI222 U1593 ( .A(n3218), .B(n6501), .C(n6320), .D(n3219), .Q(n3217) );
  OAI222 U1595 ( .A(n4929), .B(n6585), .C(n4928), .D(n6582), .Q(n3223) );
  OAI222 U1596 ( .A(n5223), .B(n6575), .C(n5222), .D(n6573), .Q(n3222) );
  OAI222 U1597 ( .A(n5225), .B(n6566), .C(n5224), .D(n6563), .Q(n3221) );
  OAI222 U1598 ( .A(n5227), .B(n6557), .C(n5226), .D(n6554), .Q(n3220) );
  OAI222 U1600 ( .A(n4881), .B(n6585), .C(n4880), .D(n6581), .Q(n3227) );
  OAI222 U1601 ( .A(n5069), .B(n6575), .C(n5068), .D(n6572), .Q(n3226) );
  OAI222 U1603 ( .A(n5073), .B(n6557), .C(n5072), .D(n6554), .Q(n3224) );
  OAI222 U1604 ( .A(n4681), .B(n6418), .C(n4680), .D(n6420), .Q(n3216) );
  OAI222 U1605 ( .A(n4679), .B(n6414), .C(n4678), .D(n6416), .Q(n3215) );
  OAI212 U1606 ( .A(n6402), .B(n5953), .C(n3228), .Q(n3214) );
  OAI222 U1609 ( .A(n1170), .B(n6005), .C(n6401), .D(n5881), .Q(n3230) );
  OAI222 U1610 ( .A(n4786), .B(n6392), .C(n6398), .D(n5980), .Q(n3229) );
  OAI222 U1615 ( .A(n3239), .B(n6501), .C(n6319), .D(n3240), .Q(n3238) );
  OAI222 U1617 ( .A(n4943), .B(n6585), .C(n4942), .D(n6581), .Q(n3244) );
  OAI222 U1618 ( .A(n5265), .B(n6575), .C(n5264), .D(n6572), .Q(n3243) );
  OAI222 U1619 ( .A(n5267), .B(n6566), .C(n5266), .D(n6563), .Q(n3242) );
  OAI222 U1620 ( .A(n5269), .B(n6557), .C(n5268), .D(n6554), .Q(n3241) );
  OAI222 U1622 ( .A(n4903), .B(n6585), .C(n4902), .D(n6581), .Q(n3248) );
  OAI222 U1623 ( .A(n5139), .B(n6575), .C(n5138), .D(n6572), .Q(n3247) );
  OAI222 U1624 ( .A(n5141), .B(n6566), .C(n5140), .D(n6564), .Q(n3246) );
  OAI222 U1625 ( .A(n5143), .B(n6557), .C(n5142), .D(n6555), .Q(n3245) );
  OAI222 U1626 ( .A(n4685), .B(n1937), .C(n4684), .D(n1938), .Q(n3237) );
  OAI222 U1627 ( .A(n4683), .B(n1939), .C(n4682), .D(n1940), .Q(n3236) );
  OAI212 U1628 ( .A(n1941), .B(n5952), .C(n3249), .Q(n3235) );
  OAI222 U1631 ( .A(n1170), .B(n6004), .C(n6400), .D(n5880), .Q(n3251) );
  OAI222 U1632 ( .A(n4814), .B(n1949), .C(n6398), .D(n5979), .Q(n3250) );
  OAI222 U1637 ( .A(n3260), .B(n6501), .C(n6319), .D(n3261), .Q(n3259) );
  OAI222 U1639 ( .A(n4885), .B(n6585), .C(n4884), .D(n6581), .Q(n3265) );
  OAI222 U1640 ( .A(n5081), .B(n6575), .C(n5080), .D(n6572), .Q(n3264) );
  OAI222 U1641 ( .A(n5083), .B(n6566), .C(n5082), .D(n1930), .Q(n3263) );
  OAI222 U1642 ( .A(n5085), .B(n6557), .C(n5084), .D(n6554), .Q(n3262) );
  OAI222 U1644 ( .A(n5347), .B(n6584), .C(n5346), .D(n6581), .Q(n3269) );
  OAI222 U1645 ( .A(n4969), .B(n6574), .C(n4968), .D(n6572), .Q(n3268) );
  OAI222 U1648 ( .A(n4689), .B(n6419), .C(n4688), .D(n6421), .Q(n3258) );
  OAI222 U1649 ( .A(n4687), .B(n6415), .C(n4686), .D(n6417), .Q(n3257) );
  OAI212 U1650 ( .A(n6403), .B(n5951), .C(n3270), .Q(n3256) );
  OAI222 U1653 ( .A(n1170), .B(n6003), .C(n1948), .D(n5879), .Q(n3272) );
  OAI222 U1654 ( .A(n4722), .B(n6393), .C(n6396), .D(n5978), .Q(n3271) );
  OAI222 U1659 ( .A(n3281), .B(n6501), .C(n6319), .D(n3282), .Q(n3280) );
  OAI222 U1661 ( .A(n4923), .B(n6584), .C(n4922), .D(n6581), .Q(n3286) );
  OAI222 U1662 ( .A(n5207), .B(n6574), .C(n5206), .D(n6572), .Q(n3285) );
  OAI222 U1663 ( .A(n5209), .B(n6565), .C(n5208), .D(n1930), .Q(n3284) );
  OAI222 U1664 ( .A(n5211), .B(n6556), .C(n5210), .D(n6555), .Q(n3283) );
  OAI222 U1666 ( .A(n4875), .B(n6584), .C(n4874), .D(n6581), .Q(n3290) );
  OAI222 U1667 ( .A(n5051), .B(n6574), .C(n5050), .D(n6572), .Q(n3289) );
  OAI222 U1669 ( .A(n5055), .B(n6556), .C(n5054), .D(n6555), .Q(n3287) );
  OAI222 U1670 ( .A(n4697), .B(n6418), .C(n4696), .D(n6420), .Q(n3279) );
  OAI222 U1671 ( .A(n4695), .B(n6414), .C(n4694), .D(n6416), .Q(n3278) );
  OAI212 U1672 ( .A(n6402), .B(n5950), .C(n3291), .Q(n3277) );
  OAI222 U1675 ( .A(n1170), .B(n6002), .C(n6401), .D(n5878), .Q(n3293) );
  OAI222 U1676 ( .A(n4778), .B(n6392), .C(n6398), .D(n5977), .Q(n3292) );
  OAI222 U1681 ( .A(n3302), .B(n6501), .C(n6319), .D(n3303), .Q(n3301) );
  OAI222 U1683 ( .A(n4937), .B(n6584), .C(n4936), .D(n6581), .Q(n3307) );
  OAI222 U1684 ( .A(n5247), .B(n6574), .C(n5246), .D(n6572), .Q(n3306) );
  OAI222 U1685 ( .A(n5249), .B(n6565), .C(n5248), .D(n1930), .Q(n3305) );
  OAI222 U1686 ( .A(n5251), .B(n6556), .C(n5250), .D(n6554), .Q(n3304) );
  OAI222 U1688 ( .A(n4893), .B(n6584), .C(n4892), .D(n6581), .Q(n3311) );
  OAI222 U1689 ( .A(n5111), .B(n6574), .C(n5110), .D(n6572), .Q(n3310) );
  OAI222 U1690 ( .A(n5113), .B(n6565), .C(n5112), .D(n6564), .Q(n3309) );
  OAI222 U1691 ( .A(n5115), .B(n6556), .C(n5114), .D(n6555), .Q(n3308) );
  OAI222 U1692 ( .A(n4701), .B(n1937), .C(n4700), .D(n1938), .Q(n3300) );
  OAI222 U1693 ( .A(n4699), .B(n1939), .C(n4698), .D(n1940), .Q(n3299) );
  OAI212 U1694 ( .A(n1941), .B(n5949), .C(n3312), .Q(n3298) );
  OAI222 U1697 ( .A(n1170), .B(n6001), .C(n6400), .D(n5877), .Q(n3314) );
  OAI222 U1698 ( .A(n4802), .B(n1949), .C(n6398), .D(n5976), .Q(n3313) );
  OAI222 U1703 ( .A(n3323), .B(n6501), .C(n6319), .D(n3324), .Q(n3322) );
  OAI222 U1705 ( .A(n4905), .B(n6584), .C(n4904), .D(n6581), .Q(n3328) );
  OAI222 U1706 ( .A(n5145), .B(n6574), .C(n5144), .D(n6572), .Q(n3327) );
  OAI222 U1707 ( .A(n5147), .B(n6565), .C(n5146), .D(n1930), .Q(n3326) );
  OAI222 U1708 ( .A(n5149), .B(n6556), .C(n5148), .D(n6555), .Q(n3325) );
  OAI222 U1710 ( .A(n4855), .B(n6584), .C(n4854), .D(n6581), .Q(n3332) );
  OAI222 U1711 ( .A(n4997), .B(n6574), .C(n4996), .D(n6572), .Q(n3331) );
  OAI222 U1712 ( .A(n4999), .B(n6565), .C(n4998), .D(n1930), .Q(n3330) );
  OAI222 U1713 ( .A(n5349), .B(n6556), .C(n5348), .D(n6554), .Q(n3329) );
  OAI222 U1714 ( .A(n4705), .B(n6419), .C(n4704), .D(n6421), .Q(n3321) );
  OAI222 U1715 ( .A(n4703), .B(n6415), .C(n4702), .D(n6417), .Q(n3320) );
  OAI212 U1716 ( .A(n1941), .B(n5948), .C(n3333), .Q(n3319) );
  OAI222 U1719 ( .A(n1170), .B(n6000), .C(n1948), .D(n5876), .Q(n3335) );
  OAI222 U1720 ( .A(n4742), .B(n6393), .C(n6397), .D(n5975), .Q(n3334) );
  OAI222 U1725 ( .A(n3344), .B(n6498), .C(n6319), .D(n3345), .Q(n3343) );
  OAI222 U1727 ( .A(n5331), .B(n6584), .C(n5330), .D(n6581), .Q(n3349) );
  OAI222 U1728 ( .A(n5287), .B(n6574), .C(n5286), .D(n6572), .Q(n3348) );
  OAI222 U1729 ( .A(n5289), .B(n6565), .C(n5288), .D(n6564), .Q(n3347) );
  OAI222 U1730 ( .A(n5291), .B(n6556), .C(n5290), .D(n6554), .Q(n3346) );
  OAI222 U1732 ( .A(n4837), .B(n6584), .C(n4836), .D(n6581), .Q(n3353) );
  OAI222 U1735 ( .A(n4949), .B(n6574), .C(n4948), .D(n6572), .Q(n3352) );
  OAI222 U1738 ( .A(n4951), .B(n6565), .C(n4950), .D(n1930), .Q(n3351) );
  OAI222 U1742 ( .A(n5315), .B(n6556), .C(n5314), .D(n6555), .Q(n3350) );
  OAI222 U1746 ( .A(n4709), .B(n6418), .C(n4708), .D(n6420), .Q(n3342) );
  OAI222 U1749 ( .A(n4707), .B(n6414), .C(n4706), .D(n6416), .Q(n3341) );
  OAI212 U1752 ( .A(n6402), .B(n5947), .C(n3363), .Q(n3340) );
  OAI222 U1758 ( .A(n1170), .B(n5898), .C(n5692), .D(n6400), .Q(n3367) );
  OAI222 U1762 ( .A(n4830), .B(n6392), .C(n6396), .D(n5974), .Q(n3366) );
  OAI212 U1785 ( .A(n3374), .B(n3375), .C(n6084), .Q(
        \instruction_decode/hazard_unit/n5 ) );
  OAI222 U1810 ( .A(n3407), .B(n3408), .C(n3409), .D(n3410), .Q(n3406) );
  OAI222 U1812 ( .A(n1285), .B(n3414), .C(n1284), .D(n1326), .Q(n3413) );
  OAI212 U1816 ( .A(n3419), .B(n3398), .C(n3420), .Q(n3418) );
  OAI212 U1817 ( .A(n6514), .B(n3421), .C(n3422), .Q(n3405) );
  OAI222 U1832 ( .A(n3448), .B(n3410), .C(n6514), .D(n3449), .Q(n3447) );
  OAI222 U1834 ( .A(n1263), .B(n3415), .C(n1264), .D(n3414), .Q(n3452) );
  OAI222 U1835 ( .A(n1268), .B(n1326), .C(n1269), .D(n1322), .Q(n3451) );
  OAI212 U1840 ( .A(n1253), .B(n3445), .C(n3463), .Q(n3461) );
  XOR31 U1846 ( .A(n3471), .B(n1360), .C(n3472), .Q(n3470) );
  OAI212 U1865 ( .A(n6514), .B(n6348), .C(n1301), .Q(n3506) );
  OAI222 U1877 ( .A(n1356), .B(n6352), .C(n3526), .D(n3407), .Q(n3525) );
  XOR31 U1878 ( .A(n3515), .B(n1356), .C(n3516), .Q(n3526) );
  OAI222 U1883 ( .A(n1287), .B(n3534), .C(n1251), .D(n3535), .Q(n3524) );
  OAI222 U1894 ( .A(n1263), .B(n3540), .C(n1344), .D(n3555), .Q(n3551) );
  OAI222 U1897 ( .A(n3558), .B(n3407), .C(n1420), .D(n3559), .Q(n3550) );
  OAI222 U1904 ( .A(n3569), .B(n1856), .C(n1261), .D(n3570), .Q(n3568) );
  OAI222 U1906 ( .A(n1233), .B(n3445), .C(n1228), .D(n3390), .Q(n3567) );
  OAI222 U1911 ( .A(n1275), .B(n3554), .C(n1277), .D(n3540), .Q(n3582) );
  XOR31 U1914 ( .A(n3587), .B(n1338), .C(n3588), .Q(n3586) );
  OAI222 U1926 ( .A(n1244), .B(n3604), .C(n1242), .D(n3605), .Q(n3597) );
  OAI212 U1930 ( .A(n3608), .B(n3609), .C(n1321), .Q(n3577) );
  OAI222 U1931 ( .A(n1420), .B(n3610), .C(n1418), .D(n3611), .Q(n3609) );
  OAI222 U1940 ( .A(n1461), .B(n6515), .C(n3402), .D(n3622), .Q(n3621) );
  OAI222 U1941 ( .A(n3623), .B(n3407), .C(n3624), .D(n3445), .Q(n1993) );
  XOR31 U1942 ( .A(n3625), .B(n3626), .C(n6351), .Q(n3623) );
  AOI2112 U1943 ( .A(n3628), .B(n1412), .C(n3629), .D(n3630), .Q(n3626) );
  OAI212 U1946 ( .A(n3637), .B(n3632), .C(n3638), .Q(n3636) );
  OAI212 U1953 ( .A(\execute/alu/sll_175/ML_int[3][23] ), .B(n6756), .C(n3648), 
        .Q(n3647) );
  OAI222 U1955 ( .A(\execute/alu/sll_175/ML_int[2][27] ), .B(n6759), .C(
        \execute/alu/sll_175/ML_int[2][31] ), .D(n6758), .Q(n3649) );
  OAI222 U1961 ( .A(n1307), .B(n1412), .C(n3660), .D(n3661), .Q(n3654) );
  OAI212 U1971 ( .A(n1410), .B(n3670), .C(n3671), .Q(n3669) );
  OAI212 U1985 ( .A(n1309), .B(n3689), .C(n3690), .Q(n3590) );
  OAI212 U1990 ( .A(n3697), .B(n3698), .C(n1321), .Q(n3696) );
  OAI222 U1997 ( .A(n1237), .B(n3604), .C(n1235), .D(n3605), .Q(n3699) );
  OAI222 U2008 ( .A(n3715), .B(n3716), .C(n1458), .D(n3717), .Q(n3714) );
  OAI212 U2015 ( .A(n3670), .B(n1410), .C(n3668), .Q(n3723) );
  OAI212 U2019 ( .A(n3724), .B(n3725), .C(n3672), .Q(n3671) );
  OAI222 U2024 ( .A(n1457), .B(n3733), .C(n3407), .D(n3734), .Q(n3732) );
  OAI212 U2027 ( .A(n1408), .B(n3737), .C(n3738), .Q(n3725) );
  OAI212 U2031 ( .A(n1409), .B(n3726), .C(n3672), .Q(n3735) );
  OAI222 U2042 ( .A(n3754), .B(n3755), .C(n1456), .D(n3756), .Q(n3753) );
  OAI212 U2056 ( .A(n1346), .B(n3765), .C(n3766), .Q(n3674) );
  OAI212 U2065 ( .A(n3782), .B(n6512), .C(n1454), .Q(n3768) );
  OAI222 U2068 ( .A(n3778), .B(n3741), .C(n1304), .D(n3785), .Q(n3784) );
  OAI222 U2077 ( .A(n3792), .B(n3793), .C(n1453), .D(n3794), .Q(n3791) );
  OAI212 U2087 ( .A(n3804), .B(n1400), .C(n1399), .Q(n3803) );
  OAI212 U2096 ( .A(n6199), .B(n3617), .C(n3813), .Q(n3812) );
  OAI212 U2109 ( .A(n1397), .B(n3826), .C(n3804), .Q(n3823) );
  OAI222 U2112 ( .A(n1401), .B(n3404), .C(n3811), .D(n6358), .Q(n3820) );
  OAI212 U2115 ( .A(n1340), .B(n1346), .C(n3766), .Q(n3772) );
  OAI212 U2116 ( .A(n3465), .B(n3617), .C(n3835), .Q(n3833) );
  OAI212 U2118 ( .A(n1245), .B(n3601), .C(n3836), .Q(n3486) );
  OAI222 U2125 ( .A(n1398), .B(n6514), .C(n3832), .D(n6358), .Q(n3842) );
  OAI212 U2132 ( .A(n1398), .B(n3827), .C(n3640), .Q(n3844) );
  OAI222 U2136 ( .A(n1396), .B(n6352), .C(n6348), .D(n3617), .Q(n3856) );
  OAI212 U2137 ( .A(n3407), .B(n3857), .C(n3858), .Q(n3855) );
  OAI212 U2139 ( .A(n1238), .B(n3601), .C(n3860), .Q(n3498) );
  OAI212 U2148 ( .A(n3872), .B(n3873), .C(n3874), .Q(n3848) );
  OAI212 U2150 ( .A(n3876), .B(n3870), .C(n3877), .Q(n3854) );
  OAI212 U2154 ( .A(n1450), .B(n3880), .C(n3881), .Q(n3853) );
  OAI212 U2167 ( .A(n1257), .B(n3605), .C(n3896), .Q(n3533) );
  OAI222 U2179 ( .A(n1265), .B(n1346), .C(n3407), .D(n3908), .Q(n3905) );
  OAI212 U2195 ( .A(n1230), .B(n3601), .C(n3920), .Q(n3572) );
  OAI212 U2199 ( .A(n1246), .B(n3390), .C(n3927), .Q(n3926) );
  OAI212 U2200 ( .A(n3928), .B(n3929), .C(n1321), .Q(n3927) );
  OAI222 U2202 ( .A(n1418), .B(n6508), .C(n1420), .D(n6511), .Q(n3928) );
  OAI212 U2203 ( .A(n1310), .B(n6352), .C(n3932), .Q(n3925) );
  OAI212 U2224 ( .A(n1310), .B(n6517), .C(n3438), .Q(n3952) );
  OAI212 U2236 ( .A(n1447), .B(n3965), .C(n3766), .Q(n3964) );
  OAI222 U2238 ( .A(n1279), .B(n1346), .C(n3407), .D(n3967), .Q(n3963) );
  OAI212 U2259 ( .A(n3407), .B(n3988), .C(n3989), .Q(n3986) );
  OAI212 U2271 ( .A(n1382), .B(n4000), .C(n3975), .Q(n3996) );
  OAI212 U2272 ( .A(n4001), .B(n4002), .C(n4003), .Q(n3975) );
  OAI212 U2273 ( .A(n4004), .B(n3999), .C(n4005), .Q(n3985) );
  OAI212 U2279 ( .A(n1445), .B(n4008), .C(n4009), .Q(n3984) );
  OAI212 U2313 ( .A(n4039), .B(n6514), .C(n4042), .Q(n4034) );
  AOI2112 U2316 ( .A(n4044), .B(n4045), .C(n4046), .D(n4047), .Q(n4041) );
  AOI212 U2319 ( .A(n4053), .B(n4054), .C(n4055), .Q(n4051) );
  OAI222 U2333 ( .A(n1278), .B(n3540), .C(n3407), .D(n4076), .Q(n4074) );
  OAI222 U2340 ( .A(n1439), .B(n4081), .C(n3624), .D(n4082), .Q(n4073) );
  OAI212 U2344 ( .A(n4085), .B(n4086), .C(n1473), .Q(n3766) );
  OAI222 U2347 ( .A(n1377), .B(n6352), .C(n6514), .D(n4091), .Q(n4090) );
  OAI222 U2354 ( .A(n1271), .B(n3534), .C(n1239), .D(n3535), .Q(n4098) );
  OAI212 U2358 ( .A(n3995), .B(n4105), .C(n4106), .Q(n4104) );
  OAI222 U2360 ( .A(n1436), .B(n4107), .C(n3407), .D(n4108), .Q(n4103) );
  OAI222 U2373 ( .A(n1285), .B(n3554), .C(n1286), .D(n3540), .Q(n4120) );
  OAI212 U2380 ( .A(n1257), .B(n4082), .C(n4125), .Q(n4119) );
  OAI212 U2381 ( .A(n4126), .B(n4127), .C(n4128), .Q(n4125) );
  OAI222 U2382 ( .A(n6346), .B(n3404), .C(n1434), .D(n6517), .Q(n4127) );
  OAI212 U2384 ( .A(n3659), .B(n4131), .C(n4132), .Q(n3713) );
  OAI222 U2386 ( .A(n1288), .B(n4105), .C(n1434), .D(n4133), .Q(n4118) );
  OAI212 U2388 ( .A(n5821), .B(n3622), .C(n4135), .Q(n3720) );
  OAI222 U2390 ( .A(n4136), .B(n3407), .C(n6358), .D(n4137), .Q(n4117) );
  OAI222 U2399 ( .A(n1284), .B(n3570), .C(n1250), .D(n3445), .Q(n4141) );
  OAI222 U2422 ( .A(n1264), .B(n3554), .C(n1266), .D(n3540), .Q(n4161) );
  OAI222 U2423 ( .A(n1370), .B(n4162), .C(n1227), .D(n4082), .Q(n4160) );
  OAI222 U2426 ( .A(n6345), .B(n3404), .C(n6210), .D(n6517), .Q(n4164) );
  OAI222 U2428 ( .A(n1267), .B(n4105), .C(n6210), .D(n4166), .Q(n4159) );
  OAI222 U2430 ( .A(n4167), .B(n3407), .C(n6358), .D(n4168), .Q(n4158) );
  AOI2112 U2434 ( .A(n4170), .B(n4171), .C(n4172), .D(n4173), .Q(n4063) );
  AOI212 U2435 ( .A(n3443), .B(n3420), .C(n4174), .Q(n4173) );
  OAI222 U2437 ( .A(n3419), .B(n3398), .C(n4175), .D(n4176), .Q(n4174) );
  OAI222 U2462 ( .A(n1280), .B(n3540), .C(n1430), .D(n4196), .Q(n4184) );
  OAI222 U2468 ( .A(n1278), .B(n4105), .C(n6344), .D(n4200), .Q(n4183) );
  OAI212 U2499 ( .A(n3553), .B(n3765), .C(n3504), .Q(n4102) );
  OAI212 U2503 ( .A(n1239), .B(n3431), .C(n4224), .Q(n4223) );
  OAI212 U2511 ( .A(n4232), .B(n4233), .C(n1366), .Q(n4231) );
  OAI212 U2517 ( .A(n1297), .B(n4235), .C(n3420), .Q(n4216) );
  OAI212 U2521 ( .A(n3442), .B(n3440), .C(n3443), .Q(n4237) );
  OAI212 U2524 ( .A(n3471), .B(n6250), .C(n4239), .Q(n4050) );
  AOI222 U2525 ( .A(n4240), .B(n4241), .C(n4242), .D(n3467), .Q(n4239) );
  AOI212 U2533 ( .A(n3471), .B(n1360), .C(n4243), .Q(n4240) );
  OAI2112 U2539 ( .A(n3938), .B(n6341), .C(n6321), .D(n1311), .Q(n4053) );
  OAI2112 U2542 ( .A(n6204), .B(n3692), .C(n3589), .D(n4247), .Q(n4244) );
  XNR22 U2550 ( .A(n3627), .B(n6349), .Q(n3587) );
  OAI222 U2577 ( .A(n3995), .B(n3417), .C(n3416), .D(n1274), .Q(n4262) );
  OAI222 U2583 ( .A(n1460), .B(n3611), .C(n1461), .D(n1293), .Q(n3995) );
  OAI212 U2610 ( .A(n3718), .B(n3716), .C(n4292), .Q(n4284) );
  OAI212 U2611 ( .A(n1457), .B(n1409), .C(n4293), .Q(n4292) );
  OAI212 U2613 ( .A(n1454), .B(n1405), .C(n4296), .Q(n4295) );
  OAI222 U2622 ( .A(n4313), .B(n4314), .C(n4315), .D(n1373), .Q(n4312) );
  OAI212 U2624 ( .A(n6346), .B(n1372), .C(n4316), .Q(n4314) );
  OAI212 U2628 ( .A(n6345), .B(n1370), .C(n4317), .Q(n4313) );
  OAI222 U2649 ( .A(n1428), .B(n1366), .C(n6344), .D(n1367), .Q(n4318) );
  OAI222 U2650 ( .A(n6210), .B(n4338), .C(n1430), .D(n4170), .Q(n4323) );
  OAI212 U2651 ( .A(n1439), .B(n4083), .C(n1384), .Q(n4311) );
  OAI222 U2652 ( .A(n1445), .B(n1385), .C(n4340), .D(n4339), .Q(n4309) );
  OAI222 U2656 ( .A(n3907), .B(n3911), .C(n3966), .D(n3972), .Q(n4306) );
  OAI222 U2666 ( .A(n4333), .B(n4341), .C(n1414), .D(n4342), .Q(n4278) );
  OAI212 U2670 ( .A(n1259), .B(n6517), .C(n3438), .Q(n4344) );
  OAI212 U2672 ( .A(n1262), .B(n3553), .C(n4345), .Q(n4277) );
  OAI222 U2710 ( .A(n1233), .B(n4372), .C(n1234), .D(n3604), .Q(n4368) );
  OAI212 U2759 ( .A(n4398), .B(n4399), .C(n1321), .Q(n4382) );
  OAI212 U2796 ( .A(n4409), .B(n5946), .C(n6247), .Q(n4414) );
  OAI222 U2806 ( .A(n5696), .B(n6489), .C(n1419), .D(n5942), .Q(\execute/n459 ) );
  AOI222 U2810 ( .A(n6075), .B(n6490), .C(\execute/op_21 [9]), .D(n6489), .Q(
        n4236) );
  OAI212 U2811 ( .A(n6950), .B(n5832), .C(n4426), .Q(\execute/op_21 [9]) );
  AOI222 U2813 ( .A(n6074), .B(n6490), .C(\execute/op_21 [8]), .D(n5734), .Q(
        n3439) );
  OAI212 U2814 ( .A(n6948), .B(n5832), .C(n4429), .Q(\execute/op_21 [8]) );
  OAI212 U2817 ( .A(n6946), .B(n5832), .C(n4430), .Q(\execute/op_21 [7]) );
  OAI212 U2820 ( .A(n6944), .B(n5831), .C(n4431), .Q(\execute/op_21 [6]) );
  AOI222 U2822 ( .A(n6246), .B(n6490), .C(\execute/op_21 [5]), .D(n6489), .Q(
        n3538) );
  OAI212 U2823 ( .A(n6942), .B(n5832), .C(n4432), .Q(\execute/op_21 [5]) );
  AOI222 U2824 ( .A(n6333), .B(data_2[5]), .C(n5815), .D(ram_adr[5]), .Q(n4432) );
  OAI222 U2825 ( .A(n6927), .B(n5638), .C(n5828), .D(n5639), .Q(
        write_data_reg[5]) );
  OAI222 U2826 ( .A(n5695), .B(n6489), .C(n1421), .D(n5942), .Q(\execute/n453 ) );
  OAI212 U2827 ( .A(n6940), .B(n5832), .C(n4433), .Q(\execute/op_21 [4]) );
  OAI212 U2830 ( .A(n6992), .B(n5832), .C(n4434), .Q(\execute/op_21 [30]) );
  AOI222 U2832 ( .A(n6232), .B(n6490), .C(\execute/op_21 [2]), .D(n6489), .Q(
        n3681) );
  OAI212 U2833 ( .A(n6935), .B(n5831), .C(n4435), .Q(\execute/op_21 [2]) );
  OAI212 U2836 ( .A(n6990), .B(n5832), .C(n4436), .Q(\execute/op_21 [29]) );
  OAI212 U2839 ( .A(n6988), .B(n5832), .C(n4437), .Q(\execute/op_21 [28]) );
  OAI212 U2842 ( .A(n6986), .B(n5832), .C(n4438), .Q(\execute/op_21 [27]) );
  OAI212 U2845 ( .A(n6984), .B(n5832), .C(n4439), .Q(\execute/op_21 [26]) );
  OAI212 U2848 ( .A(n6982), .B(n5832), .C(n4440), .Q(\execute/op_21 [25]) );
  OAI212 U2851 ( .A(n6980), .B(n5832), .C(n4441), .Q(\execute/op_21 [24]) );
  OAI212 U2854 ( .A(n6978), .B(n5832), .C(n4442), .Q(\execute/op_21 [23]) );
  OAI212 U2857 ( .A(n6976), .B(n5832), .C(n4443), .Q(\execute/op_21 [22]) );
  OAI212 U2860 ( .A(n6974), .B(n5831), .C(n4445), .Q(\execute/op_21 [21]) );
  OAI212 U2863 ( .A(n6972), .B(n5832), .C(n4446), .Q(\execute/op_21 [20]) );
  AOI222 U2865 ( .A(n6247), .B(n6490), .C(\execute/op_21 [1]), .D(n6489), .Q(
        n3930) );
  OAI212 U2866 ( .A(n6933), .B(n5831), .C(n4447), .Q(\execute/op_21 [1]) );
  OAI212 U2869 ( .A(n6970), .B(n4425), .C(n4448), .Q(\execute/op_21 [19]) );
  OAI212 U2872 ( .A(n6968), .B(n5832), .C(n4449), .Q(\execute/op_21 [18]) );
  OAI212 U2875 ( .A(n6966), .B(n5832), .C(n4450), .Q(\execute/op_21 [17]) );
  OAI212 U2878 ( .A(n6964), .B(n5832), .C(n4451), .Q(\execute/op_21 [16]) );
  OAI222 U2880 ( .A(n5619), .B(n6489), .C(n1440), .D(n6490), .Q(\execute/n434 ) );
  OAI212 U2881 ( .A(n6962), .B(n5831), .C(n4452), .Q(\execute/op_21 [15]) );
  OAI222 U2883 ( .A(n5609), .B(n6489), .C(n1437), .D(n5942), .Q(\execute/n433 ) );
  OAI212 U2884 ( .A(n6960), .B(n5831), .C(n4453), .Q(\execute/op_21 [14]) );
  OAI222 U2886 ( .A(n5610), .B(n6489), .C(n1435), .D(n5942), .Q(\execute/n432 ) );
  OAI212 U2887 ( .A(n6958), .B(n5832), .C(n4454), .Q(\execute/op_21 [13]) );
  OAI222 U2889 ( .A(n5620), .B(n6489), .C(n1433), .D(n5942), .Q(\execute/n431 ) );
  OAI212 U2890 ( .A(n6956), .B(n5832), .C(n4455), .Q(\execute/op_21 [12]) );
  OAI222 U2892 ( .A(n5617), .B(n6489), .C(n1431), .D(n5942), .Q(\execute/n430 ) );
  OAI212 U2893 ( .A(n6954), .B(n5832), .C(n4456), .Q(\execute/op_21 [11]) );
  AOI222 U2895 ( .A(n6073), .B(n6490), .C(\execute/op_21 [10]), .D(n6489), .Q(
        n4227) );
  OAI212 U2896 ( .A(n6952), .B(n5831), .C(n4457), .Q(\execute/op_21 [10]) );
  OAI2112 U2905 ( .A(n6938), .B(n6505), .C(n4461), .D(n4462), .Q(n3592) );
  AOI222 U2907 ( .A(ram_adr[3]), .B(n6337), .C(n6340), .D(data_1[3]), .Q(n4461) );
  OAI222 U2908 ( .A(n6926), .B(n5648), .C(n5828), .D(n5649), .Q(
        write_data_reg[3]) );
  OAI2112 U2914 ( .A(n6935), .B(n6505), .C(n4465), .D(n4466), .Q(n3683) );
  OAI2112 U2921 ( .A(n6933), .B(n6505), .C(n4467), .D(n4468), .Q(n3692) );
  OAI212 U2926 ( .A(n4458), .B(n1259), .C(n4401), .Q(
        \execute/alu/sll_175/temp_int_SH[0] ) );
  OAI222 U2946 ( .A(n6926), .B(n5684), .C(n5828), .D(n5685), .Q(
        write_data_reg[11]) );
  OAI222 U2950 ( .A(n6926), .B(n5676), .C(n6924), .D(n5677), .Q(
        write_data_reg[12]) );
  OAI222 U2954 ( .A(n6926), .B(n5660), .C(n6924), .D(n5661), .Q(
        write_data_reg[20]) );
  OAI222 U2959 ( .A(n6926), .B(n5664), .C(n6924), .D(n5665), .Q(
        write_data_reg[14]) );
  OAI222 U2963 ( .A(n6926), .B(n5668), .C(n6924), .D(n5669), .Q(
        write_data_reg[15]) );
  OAI222 U2967 ( .A(n6926), .B(n5686), .C(n6924), .D(n5687), .Q(
        write_data_reg[13]) );
  OAI222 U2971 ( .A(n6926), .B(n5680), .C(n6924), .D(n5681), .Q(
        write_data_reg[10]) );
  OAI222 U2976 ( .A(n6927), .B(n5670), .C(n6924), .D(n5671), .Q(
        write_data_reg[19]) );
  OAI222 U2980 ( .A(n6927), .B(n5646), .C(n6924), .D(n5647), .Q(
        write_data_reg[21]) );
  OAI222 U2984 ( .A(n6927), .B(n5678), .C(n6924), .D(n5679), .Q(
        write_data_reg[16]) );
  OAI222 U2989 ( .A(n6927), .B(n5636), .C(n6924), .D(n5637), .Q(
        write_data_reg[26]) );
  OAI222 U2993 ( .A(n6927), .B(n5654), .C(n6924), .D(n5655), .Q(
        write_data_reg[18]) );
  OAI222 U2997 ( .A(n6927), .B(n5682), .C(n6924), .D(n5683), .Q(
        write_data_reg[17]) );
  OAI222 U3002 ( .A(n6927), .B(n5650), .C(n6924), .D(n5651), .Q(
        write_data_reg[23]) );
  OAI222 U3006 ( .A(n6927), .B(n5656), .C(n6923), .D(n5657), .Q(
        write_data_reg[24]) );
  OAI222 U3010 ( .A(n6927), .B(n5688), .C(n6923), .D(n5689), .Q(
        write_data_reg[6]) );
  OAI222 U3015 ( .A(n6927), .B(n5652), .C(n6923), .D(n5653), .Q(
        write_data_reg[22]) );
  OAI222 U3019 ( .A(n6927), .B(n5632), .C(n6923), .D(n5633), .Q(
        write_data_reg[27]) );
  OAI222 U3023 ( .A(n6928), .B(n5662), .C(n6923), .D(n5663), .Q(
        write_data_reg[25]) );
  OAI222 U3032 ( .A(n6928), .B(n5628), .C(n6923), .D(n5629), .Q(
        write_data_reg[28]) );
  OAI222 U3036 ( .A(n6928), .B(n5630), .C(n6923), .D(n5631), .Q(
        write_data_reg[29]) );
  OAI222 U3041 ( .A(n5674), .B(n6928), .C(n6923), .D(n5675), .Q(
        write_data_reg[9]) );
  OAI222 U3045 ( .A(n6928), .B(n5672), .C(n6923), .D(n5673), .Q(
        write_data_reg[7]) );
  OAI222 U3049 ( .A(n6928), .B(n5666), .C(n6923), .D(n5667), .Q(
        write_data_reg[8]) );
  AOI222 U3075 ( .A(n5946), .B(n5942), .C(\execute/op_21 [0]), .D(n6489), .Q(
        n4333) );
  OAI212 U3076 ( .A(n6931), .B(n5831), .C(n4558), .Q(\execute/op_21 [0]) );
  AOI222 U3077 ( .A(n6329), .B(data_2[0]), .C(ram_adr[0]), .D(n5816), .Q(n4558) );
  OAI212 U3080 ( .A(n6994), .B(n5832), .C(n4559), .Q(\execute/op_21 [31]) );
  NOR42 U3088 ( .A(n1486), .B(n5823), .C(n4565), .D(n4564), .Q(n4563) );
  XNR22 U3095 ( .A(write_register_ex[1]), .B(n6067), .Q(n4571) );
  OAI222 U3105 ( .A(n6926), .B(n5634), .C(n6923), .D(n5635), .Q(
        write_data_reg[31]) );
  CLKIN6 U3106 ( .A(clk), .Q(n1107) );
  CLKIN6 U3418 ( .A(n5813), .Q(n1419) );
  MUX21 \execute/alu/sll_175/M1_0_2  ( .A(n1416), .B(n1415), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][2] ) );
  MUX21 \execute/alu/sll_175/M1_0_3  ( .A(n6349), .B(n1416), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][3] ) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[28]  ( .D(n6271), .E(n6762), .C(
        clk), .RN(n6610), .Q(pc_rom[28]) );
  DFE1 \instruction_fetch/inst_out_reg[2]  ( .D(n5764), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[2]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[30]  ( .D(n5801), .E(n6762), .C(
        clk), .RN(n6611), .Q(pc_rom[30]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[1]  ( .D(n5788), .E(n6762), .C(
        clk), .RN(n6611), .Q(\instruction_fetch/mux/N14 ), .QN(n4577) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[0]  ( .D(n5781), .E(n6762), .C(
        clk), .RN(n6611), .Q(\instruction_fetch/mux/N13 ), .QN(n4576) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[31]  ( .D(n6275), .E(n6762), .C(
        clk), .RN(n6611), .Q(pc_rom[31]), .QN(n4580) );
  DFE1 \instruction_fetch/inst_out_reg[13]  ( .D(n5753), .E(n6762), .C(clk), 
        .Q(inst_out[13]), .QN(n5714) );
  DFE1 \instruction_fetch/inst_out_reg[14]  ( .D(n5752), .E(n6762), .C(clk), 
        .Q(inst_out[14]), .QN(n5711) );
  DFE1 \instruction_fetch/inst_out_reg[15]  ( .D(n5751), .E(n6762), .C(clk), 
        .Q(inst_out[15]), .QN(n5710) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[29]  ( .D(n5800), .E(n6762), .C(
        clk), .RN(n6611), .Q(pc_rom[29]), .QN(n6089) );
  DFE1 \instruction_fetch/inst_out_reg[12]  ( .D(n5754), .E(n6762), .C(clk), 
        .Q(inst_out[12]), .QN(n5712) );
  DFE1 \instruction_fetch/inst_out_reg[11]  ( .D(n5755), .E(n6762), .C(clk), 
        .Q(inst_out[11]), .QN(n5713) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[24]  ( .D(n5799), .E(n6762), .C(
        clk), .RN(n6610), .Q(pc_rom[24]) );
  DFE1 \instruction_fetch/inst_out_reg[10]  ( .D(n5756), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[10]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[27]  ( .D(n5794), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6608), .Q(
        pc_rom[27]), .QN(n6090) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[25]  ( .D(n5793), .E(n6762), .C(
        clk), .RN(n6610), .Q(pc_rom[25]), .QN(n6088) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[26]  ( .D(n5786), .E(n6762), .C(
        clk), .RN(n6610), .Q(pc_rom[26]) );
  DFE1 \instruction_fetch/inst_out_reg[30]  ( .D(n5736), .E(n6762), .C(clk), 
        .QN(n5731) );
  DFE1 \instruction_fetch/inst_out_reg[9]  ( .D(n5757), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[9]) );
  DFE1 \instruction_fetch/inst_out_reg[7]  ( .D(n5759), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[7]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[20]  ( .D(n5798), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6610), .Q(
        pc_rom[20]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[22]  ( .D(n5785), .E(n6762), .C(
        clk), .RN(n6610), .Q(pc_rom[22]) );
  DFE1 \instruction_fetch/inst_out_reg[8]  ( .D(n5758), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[8]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[19]  ( .D(n5777), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6610), .Q(
        pc_rom[19]), .QN(n6082) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[21]  ( .D(n5792), .E(n6762), .C(
        clk), .RN(n6610), .Q(pc_rom[21]), .QN(n6083) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[23]  ( .D(n5779), .E(n6762), .C(
        clk), .RN(n6610), .Q(pc_rom[23]), .QN(n6087) );
  DFE1 \instruction_fetch/inst_out_reg[27]  ( .D(n5739), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(n6086), .QN(n5718)
         );
  DFE1 \instruction_fetch/inst_out_reg[29]  ( .D(n5737), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(n6085), .QN(n5717)
         );
  DFE1 \instruction_fetch/inst_out_reg[28]  ( .D(n5738), .E(n6762), .C(clk), 
        .Q(n5945), .QN(n5715) );
  DFE1 \instruction_fetch/inst_out_reg[31]  ( .D(n5735), .E(n6762), .C(clk), 
        .QN(n5730) );
  DFE1 \instruction_fetch/inst_out_reg[26]  ( .D(n5740), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(n5868), .QN(n5716)
         );
  DFE1 \instruction_fetch/inst_out_reg[5]  ( .D(n5761), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[5]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[14]  ( .D(n5791), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6609), .Q(
        pc_rom[14]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[16]  ( .D(n5784), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6609), .Q(
        pc_rom[16]) );
  DFE1 \instruction_fetch/inst_out_reg[4]  ( .D(n5762), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[4]) );
  DFE1 \instruction_fetch/inst_out_reg[6]  ( .D(n5760), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[6]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[13]  ( .D(n5775), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6609), .Q(
        pc_rom[13]), .QN(n6078) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[15]  ( .D(n5789), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6609), .Q(
        pc_rom[15]), .QN(n6079) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[17]  ( .D(n5778), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6609), .Q(
        pc_rom[17]), .QN(n6081) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[18]  ( .D(n5774), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6609), .Q(
        pc_rom[18]) );
  DFE1 \instruction_fetch/inst_out_reg[3]  ( .D(n5763), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[3]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[8]  ( .D(
        \instruction_fetch/pc_4 [8]), .E(\instruction_decode/hazard_unit/n5 ), 
        .C(clk), .RN(n6608), .Q(pc_rom[8]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[10]  ( .D(n5796), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6609), .Q(
        pc_rom[10]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[12]  ( .D(n5790), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6609), .Q(
        pc_rom[12]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[9]  ( .D(n5780), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6608), .Q(
        pc_rom[9]), .QN(n6077) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[11]  ( .D(n5795), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6609), .Q(
        pc_rom[11]), .QN(n6076) );
  DFE1 \instruction_fetch/inst_out_reg[19]  ( .D(n5747), .E(n6762), .C(clk), 
        .Q(inst_out[19]), .QN(n5722) );
  DFE1 \instruction_fetch/inst_out_reg[24]  ( .D(n5742), .E(n6762), .C(clk), 
        .Q(inst_out[24]), .QN(n5721) );
  DFE1 \instruction_fetch/inst_out_reg[16]  ( .D(n5750), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[16]), .QN(
        n5728) );
  DFE1 \instruction_fetch/inst_out_reg[17]  ( .D(n5749), .E(n6762), .C(clk), 
        .Q(inst_out[17]), .QN(n5724) );
  DFE1 \instruction_fetch/inst_out_reg[18]  ( .D(n5748), .E(n6762), .C(clk), 
        .Q(inst_out[18]), .QN(n5726) );
  DFE1 \instruction_fetch/inst_out_reg[21]  ( .D(n5745), .E(n6762), .C(clk), 
        .Q(inst_out[21]), .QN(n5725) );
  DFE1 \instruction_fetch/inst_out_reg[0]  ( .D(n5766), .E(n6762), .C(clk), 
        .Q(inst_out[0]), .QN(n5729) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[3]  ( .D(n5787), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6608), .Q(
        \instruction_fetch/n86 ), .QN(n4581) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[4]  ( .D(n5776), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6608), .Q(
        pc_rom[4]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[6]  ( .D(n5783), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6608), .Q(
        pc_rom[6]) );
  DFE1 \instruction_fetch/inst_out_reg[1]  ( .D(n5765), .E(n6762), .C(clk), 
        .Q(inst_out[1]) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[5]  ( .D(n5782), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6608), .Q(
        pc_rom[5]), .QN(n6071) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[7]  ( .D(
        \instruction_fetch/pc_4 [7]), .E(\instruction_decode/hazard_unit/n5 ), 
        .C(clk), .RN(n6608), .Q(pc_rom[7]), .QN(n6070) );
  DFEC1 \instruction_fetch/pc_REG/old_pc_reg[2]  ( .D(n5797), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .RN(n6608), .Q(
        \instruction_fetch/n87 ), .QN(n5701) );
  DFE1 \instruction_fetch/inst_out_reg[23]  ( .D(n5743), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[23]), .QN(
        n5727) );
  DFE1 \instruction_fetch/inst_out_reg[22]  ( .D(n5744), .E(n6762), .C(clk), 
        .Q(inst_out[22]), .QN(n5723) );
  DFE1 \instruction_fetch/inst_out_reg[20]  ( .D(n5746), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[20]), .QN(
        n5720) );
  DFE1 \instruction_fetch/inst_out_reg[25]  ( .D(n5741), .E(
        \instruction_decode/hazard_unit/n5 ), .C(clk), .Q(inst_out[25]), .QN(
        n5719) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][3]  ( .D(n6937), .E(
        n6847), .C(n1107), .RN(n6619), .Q(n5929) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][4]  ( .D(
        write_data_reg[4]), .E(n6846), .C(n1107), .RN(n6619), .Q(n5928) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][7]  ( .D(
        write_data_reg[7]), .E(n6846), .C(n1107), .RN(n6619), .Q(n5846) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][8]  ( .D(
        write_data_reg[8]), .E(n6846), .C(n1107), .RN(n6619), .Q(n5833) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][9]  ( .D(n6949), .E(
        n6846), .C(n1107), .RN(n6619), .Q(n5845) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][10]  ( .D(n6951), .E(
        n6846), .C(n1107), .RN(n6619), .Q(n5925) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][11]  ( .D(
        write_data_reg[11]), .E(n6845), .C(n1107), .RN(n6619), .Q(n5923) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][12]  ( .D(n6955), .E(
        n6845), .C(n1107), .RN(n6620), .Q(n5922) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][13]  ( .D(
        write_data_reg[13]), .E(n6845), .C(n1107), .RN(n6620), .Q(n5844) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][14]  ( .D(n6959), .E(
        n6845), .C(n1107), .RN(n6620), .Q(n5921) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][15]  ( .D(
        write_data_reg[15]), .E(n6845), .C(n1107), .RN(n6620), .Q(n5919) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][16]  ( .D(
        write_data_reg[16]), .E(n6845), .C(n1107), .RN(n6620), .Q(n5917) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][17]  ( .D(n6965), .E(
        n6845), .C(n1107), .RN(n6620), .Q(n5859) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][18]  ( .D(n6967), .E(
        n6844), .C(n1107), .RN(n6620), .Q(n5931) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][19]  ( .D(n6969), .E(
        n6844), .C(n1107), .RN(n6620), .Q(n6030) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][20]  ( .D(n6971), .E(
        n6844), .C(n1107), .RN(n6620), .Q(n6029) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][23]  ( .D(n6977), .E(
        n6844), .C(n1107), .RN(n6621), .Q(n5863) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][7]  ( .D(
        write_data_reg[7]), .E(n6856), .C(n1107), .RN(n6639), .Q(n5847) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][8]  ( .D(
        write_data_reg[8]), .E(n6856), .C(n1107), .RN(n6639), .Q(n5838) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][11]  ( .D(
        write_data_reg[11]), .E(n6855), .C(n1107), .RN(n6639), .Q(n5924) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][12]  ( .D(n6955), .E(
        n6855), .C(n1107), .RN(n6639), .Q(n6034) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][13]  ( .D(
        write_data_reg[13]), .E(n6855), .C(n1107), .RN(n6640), .Q(n5860) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][14]  ( .D(n6959), .E(
        n6855), .C(n1107), .RN(n6640), .Q(n6033) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][15]  ( .D(
        write_data_reg[15]), .E(n6855), .C(n1107), .RN(n6640), .Q(n5920) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][16]  ( .D(
        write_data_reg[16]), .E(n6855), .C(n1107), .RN(n6640), .Q(n5918) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][19]  ( .D(n6969), .E(
        n6854), .C(n1107), .RN(n6640), .Q(n6031) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][0]  ( .D(n6930), .E(
        n6862), .C(n1107), .RN(n6666), .Q(n5935) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][3]  ( .D(n6936), .E(
        n6862), .C(n1107), .RN(n6666), .Q(n6058) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][4]  ( .D(n6939), .E(
        n6861), .C(n1107), .RN(n6666), .Q(n6057) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][5]  ( .D(n6941), .E(
        n6861), .C(n1107), .RN(n6667), .Q(n6056) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][6]  ( .D(n6943), .E(
        n6861), .C(n1107), .RN(n6667), .Q(n6055) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][7]  ( .D(n6945), .E(
        n6861), .C(n1107), .RN(n6667), .Q(n5866) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][8]  ( .D(
        write_data_reg[8]), .E(n6861), .C(n1107), .RN(n6667), .Q(n5835) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][9]  ( .D(n6949), .E(
        n6861), .C(n1107), .RN(n6667), .Q(n5865) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][10]  ( .D(n6951), .E(
        n6861), .C(n1107), .RN(n6667), .Q(n6054) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][11]  ( .D(n6953), .E(
        n6860), .C(n1107), .RN(n6667), .Q(n6053) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][12]  ( .D(
        write_data_reg[12]), .E(n6860), .C(n1107), .RN(n6667), .Q(n6052) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][13]  ( .D(
        write_data_reg[13]), .E(n6860), .C(n1107), .RN(n6667), .Q(n5936) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][14]  ( .D(n6959), .E(
        n6860), .C(n1107), .RN(n6668), .Q(n6051) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][15]  ( .D(n6961), .E(
        n6860), .C(n1107), .RN(n6668), .Q(n6050) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][16]  ( .D(n6963), .E(
        n6860), .C(n1107), .RN(n6668), .Q(n6049) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][17]  ( .D(
        write_data_reg[17]), .E(n6860), .C(n1107), .RN(n6668), .Q(n5934) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][18]  ( .D(n6967), .E(
        n6859), .C(n1107), .RN(n6668), .Q(n6060) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][19]  ( .D(
        write_data_reg[19]), .E(n6859), .C(n1107), .RN(n6668), .Q(n5933) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][20]  ( .D(
        write_data_reg[20]), .E(n6859), .C(n1107), .RN(n6668), .Q(n5849) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][21]  ( .D(
        write_data_reg[21]), .E(n6859), .C(n1107), .RN(n6668), .Q(n5850) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][22]  ( .D(n6975), .E(
        n6859), .C(n1107), .RN(n6668), .Q(n6061) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][23]  ( .D(n6977), .E(
        n6859), .C(n1107), .RN(n6669), .Q(n5938) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][24]  ( .D(
        write_data_reg[24]), .E(n6859), .C(n1107), .RN(n6669), .Q(n5937) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][0]  ( .D(
        write_data_reg[0]), .E(n6867), .C(n1107), .RN(n6701), .Q(n6020) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][0]  ( .D(
        write_data_reg[0]), .E(n6882), .C(n1107), .RN(n6694), .QN(n5898) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][3]  ( .D(n6936), .E(
        n6882), .C(n1107), .RN(n6694), .QN(n6011) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][4]  ( .D(
        write_data_reg[4]), .E(n6881), .C(n1107), .RN(n6694), .QN(n6012) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][5]  ( .D(n6941), .E(
        n6881), .C(n1107), .RN(n6695), .QN(n6013) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][7]  ( .D(n6945), .E(
        n6881), .C(n1107), .RN(n6695), .QN(n6015) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][8]  ( .D(n6947), .E(
        n6881), .C(n1107), .RN(n6695), .QN(n6016) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][9]  ( .D(n6949), .E(
        n6881), .C(n1107), .RN(n6695), .QN(n6017) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][10]  ( .D(
        write_data_reg[10]), .E(n6881), .C(n1107), .RN(n6695), .QN(n6000) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][12]  ( .D(
        write_data_reg[12]), .E(n6880), .C(n1107), .RN(n6695), .QN(n6002) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][13]  ( .D(n6957), .E(
        n6880), .C(n1107), .RN(n6695), .QN(n6018) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][14]  ( .D(
        write_data_reg[14]), .E(n6880), .C(n1107), .RN(n6695), .QN(n6003) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][15]  ( .D(n6961), .E(
        n6880), .C(n1107), .RN(n6696), .QN(n6004) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][16]  ( .D(n6963), .E(
        n6880), .C(n1107), .RN(n6696), .QN(n6005) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][17]  ( .D(
        write_data_reg[17]), .E(n6880), .C(n1107), .RN(n6696), .QN(n5899) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][18]  ( .D(n6967), .E(
        n6880), .C(n1107), .RN(n6696), .QN(n6019) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][19]  ( .D(
        write_data_reg[19]), .E(n6879), .C(n1107), .RN(n6696), .QN(n5900) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][20]  ( .D(
        write_data_reg[20]), .E(n6879), .C(n1107), .RN(n6696), .QN(n5901) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][21]  ( .D(
        write_data_reg[21]), .E(n6879), .C(n1107), .RN(n6696), .QN(n6007) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][7]  ( .D(n6945), .E(
        n6871), .C(n1107), .RN(n6698), .QN(n5995) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][11]  ( .D(n6953), .E(
        n6870), .C(n1107), .RN(n6698), .QN(n5976) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][12]  ( .D(
        write_data_reg[12]), .E(n6870), .C(n1107), .RN(n6698), .QN(n5977) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][13]  ( .D(n6957), .E(
        n6870), .C(n1107), .RN(n6699), .QN(n5998) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][15]  ( .D(n6961), .E(
        n6870), .C(n1107), .RN(n6699), .QN(n5979) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][3]  ( .D(n6936), .E(
        n6877), .C(n1107), .RN(n6713), .QN(n5891) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][7]  ( .D(n6945), .E(
        n6876), .C(n1107), .RN(n6714), .QN(n5895) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][8]  ( .D(n6947), .E(
        n6876), .C(n1107), .RN(n6714), .QN(n5896) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][11]  ( .D(n6953), .E(
        n6875), .C(n1107), .RN(n6714), .QN(n5877) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][12]  ( .D(
        write_data_reg[12]), .E(n6875), .C(n1107), .RN(n6714), .QN(n5878) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][13]  ( .D(n6957), .E(
        n6875), .C(n1107), .RN(n6714), .QN(n5897) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][14]  ( .D(
        write_data_reg[14]), .E(n6875), .C(n1107), .RN(n6714), .QN(n5879) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][15]  ( .D(n6961), .E(
        n6875), .C(n1107), .RN(n6714), .QN(n5880) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][16]  ( .D(n6963), .E(
        n6875), .C(n1107), .RN(n6715), .QN(n5881) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][17]  ( .D(
        write_data_reg[17]), .E(n6875), .C(n1107), .RN(n6715), .QN(n5851) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][19]  ( .D(
        write_data_reg[19]), .E(n6874), .C(n1107), .RN(n6715), .QN(n5852) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][11]  ( .D(n6953), .E(
        n6878), .C(n1107), .RN(n6720), .QN(n6001) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][23]  ( .D(
        write_data_reg[23]), .E(n6878), .C(n1107), .RN(n6720), .QN(n5902) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][11]  ( .D(n6953), .E(
        n6788), .C(n1107), .RN(n6722), .QN(n5949) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][11]  ( .D(
        write_data_reg[11]), .E(n6775), .C(n1107), .RN(n6650), .QN(n4701) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][7]  ( .D(n6945), .E(
        n6851), .C(n1107), .RN(n6670), .QN(n4822) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][11]  ( .D(n6953), .E(
        n6850), .C(n1107), .RN(n6671), .QN(n4802) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][12]  ( .D(
        write_data_reg[12]), .E(n6850), .C(n1107), .RN(n6671), .QN(n4778) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][15]  ( .D(n6961), .E(
        n6850), .C(n1107), .RN(n6671), .QN(n4814) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][11]  ( .D(n6953), .E(
        n6785), .C(n1107), .RN(n6711), .Q(n5368) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][0]  ( .D(
        write_data_reg[0]), .E(n6797), .C(n1107), .RN(n6716), .Q(n5358) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][1]  ( .D(
        write_data_reg[1]), .E(n6797), .C(n1107), .RN(n6716), .Q(n5442) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][2]  ( .D(
        write_data_reg[2]), .E(n6797), .C(n1107), .RN(n6717), .Q(n5526) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][3]  ( .D(n6936), .E(n6797), .C(n1107), .RN(n6717), .Q(n5550) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][4]  ( .D(
        write_data_reg[4]), .E(n6796), .C(n1107), .RN(n6717), .Q(n5558) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][5]  ( .D(n6941), .E(n6796), .C(n1107), .RN(n6717), .Q(n5566) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][6]  ( .D(n6943), .E(n6796), .C(n1107), .RN(n6717), .Q(n5574) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][7]  ( .D(n6945), .E(n6796), .C(n1107), .RN(n6717), .Q(n5582) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][8]  ( .D(n6947), .E(n6796), .C(n1107), .RN(n6717), .Q(n5590) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][9]  ( .D(n6949), .E(n6796), .C(n1107), .RN(n6717), .Q(n5598) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][10]  ( .D(
        write_data_reg[10]), .E(n6796), .C(n1107), .RN(n6717), .Q(n5362) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][12]  ( .D(
        write_data_reg[12]), .E(n6795), .C(n1107), .RN(n6718), .Q(n5378) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][13]  ( .D(n6957), .E(
        n6795), .C(n1107), .RN(n6718), .Q(n5386) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][14]  ( .D(
        write_data_reg[14]), .E(n6795), .C(n1107), .RN(n6718), .Q(n5394) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][15]  ( .D(n6961), .E(
        n6795), .C(n1107), .RN(n6718), .Q(n5402) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][16]  ( .D(n6963), .E(
        n6795), .C(n1107), .RN(n6718), .Q(n5410) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][17]  ( .D(
        write_data_reg[17]), .E(n6795), .C(n1107), .RN(n6718), .Q(n5418) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][19]  ( .D(
        write_data_reg[19]), .E(n6794), .C(n1107), .RN(n6718), .Q(n5434) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][20]  ( .D(
        write_data_reg[20]), .E(n6794), .C(n1107), .RN(n6718), .Q(n5446) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][21]  ( .D(
        write_data_reg[21]), .E(n6794), .C(n1107), .RN(n6719), .Q(n5454) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][22]  ( .D(n6975), .E(
        n6794), .C(n1107), .RN(n6719), .Q(n5462) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][24]  ( .D(n6979), .E(
        n6794), .C(n1107), .RN(n6719), .Q(n5478) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][25]  ( .D(n6981), .E(
        n6794), .C(n1107), .RN(n6719), .Q(n5486) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][26]  ( .D(
        write_data_reg[26]), .E(n6794), .C(n1107), .RN(n6719), .Q(n5494) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][29]  ( .D(n6989), .E(
        n6793), .C(n1107), .RN(n6719), .Q(n5518) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][30]  ( .D(n6991), .E(
        n6793), .C(n1107), .RN(n6719), .Q(n5534) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][31]  ( .D(
        write_data_reg[31]), .E(n6793), .C(n1107), .RN(n6719), .Q(n5542) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][11]  ( .D(n6953), .E(
        n6793), .C(n1107), .RN(n6723), .Q(n5370) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][23]  ( .D(
        write_data_reg[23]), .E(n6793), .C(n1107), .RN(n6723), .Q(n5470) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][27]  ( .D(n6985), .E(
        n6793), .C(n1107), .RN(n6723), .Q(n5502) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][28]  ( .D(n6987), .E(
        n6793), .C(n1107), .RN(n6723), .Q(n5510) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[6][18]  ( .D(n6967), .E(
        n6795), .C(n1107), .RN(n6718), .Q(n5426) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][1]  ( .D(n6932), .E(
        n6867), .C(n1107), .RN(n6701), .Q(n5352) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][2]  ( .D(n6934), .E(
        n6867), .C(n1107), .RN(n6701), .Q(n5528) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][3]  ( .D(n6936), .E(
        n6867), .C(n1107), .RN(n6701), .Q(n5552) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][4]  ( .D(
        write_data_reg[4]), .E(n6866), .C(n1107), .RN(n6701), .Q(n5560) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][5]  ( .D(n6941), .E(
        n6866), .C(n1107), .RN(n6701), .Q(n5568) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][6]  ( .D(n6943), .E(
        n6866), .C(n1107), .RN(n6701), .Q(n5576) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][7]  ( .D(n6945), .E(
        n6866), .C(n1107), .RN(n6701), .Q(n5584) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][8]  ( .D(n6947), .E(
        n6866), .C(n1107), .RN(n6701), .Q(n5592) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][9]  ( .D(n6949), .E(
        n6866), .C(n1107), .RN(n6702), .Q(n5600) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][10]  ( .D(
        write_data_reg[10]), .E(n6866), .C(n1107), .RN(n6702), .Q(n5364) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][11]  ( .D(n6953), .E(
        n6865), .C(n1107), .RN(n6702), .Q(n5372) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][12]  ( .D(
        write_data_reg[12]), .E(n6865), .C(n1107), .RN(n6702), .Q(n5380) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][13]  ( .D(n6957), .E(
        n6865), .C(n1107), .RN(n6702), .Q(n5388) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][14]  ( .D(
        write_data_reg[14]), .E(n6865), .C(n1107), .RN(n6702), .Q(n5396) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][15]  ( .D(n6961), .E(
        n6865), .C(n1107), .RN(n6702), .Q(n5404) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][16]  ( .D(n6963), .E(
        n6865), .C(n1107), .RN(n6702), .Q(n5412) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][17]  ( .D(
        write_data_reg[17]), .E(n6865), .C(n1107), .RN(n6702), .Q(n5420) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][19]  ( .D(
        write_data_reg[19]), .E(n6864), .C(n1107), .RN(n6703), .Q(n5436) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][20]  ( .D(
        write_data_reg[20]), .E(n6864), .C(n1107), .RN(n6703), .Q(n5448) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][21]  ( .D(
        write_data_reg[21]), .E(n6864), .C(n1107), .RN(n6703), .Q(n5456) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][22]  ( .D(n6975), .E(
        n6864), .C(n1107), .RN(n6703), .Q(n5464) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][23]  ( .D(
        write_data_reg[23]), .E(n6864), .C(n1107), .RN(n6703), .Q(n5472) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][24]  ( .D(n6979), .E(
        n6864), .C(n1107), .RN(n6703), .Q(n5480) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][25]  ( .D(n6981), .E(
        n6863), .C(n1107), .RN(n6703), .Q(n5488) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][26]  ( .D(
        write_data_reg[26]), .E(n6863), .C(n1107), .RN(n6703), .Q(n5496) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][27]  ( .D(n6985), .E(
        n6863), .C(n1107), .RN(n6704), .Q(n5504) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][28]  ( .D(n6987), .E(
        n6863), .C(n1107), .RN(n6704), .Q(n5512) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][29]  ( .D(n6989), .E(
        n6863), .C(n1107), .RN(n6704), .Q(n5520) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][30]  ( .D(n6991), .E(
        n6863), .C(n1107), .RN(n6704), .Q(n5536) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][31]  ( .D(
        write_data_reg[31]), .E(n6863), .C(n1107), .RN(n6704), .Q(n5544) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[20][18]  ( .D(n6967), .E(
        n6864), .C(n1107), .RN(n6703), .Q(n5428) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][0]  ( .D(n6930), .E(
        n6847), .C(n1107), .RN(n6618), .Q(n5843) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][1]  ( .D(
        write_data_reg[1]), .E(n6847), .C(n1107), .RN(n6618), .Q(n5930) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][2]  ( .D(
        write_data_reg[2]), .E(n6847), .C(n1107), .RN(n6618), .Q(n5910) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][5]  ( .D(
        write_data_reg[5]), .E(n6846), .C(n1107), .RN(n6619), .Q(n5926) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][6]  ( .D(
        write_data_reg[6]), .E(n6846), .C(n1107), .RN(n6619), .Q(n5841) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][21]  ( .D(n6973), .E(
        n6844), .C(n1107), .RN(n6621), .Q(n5837) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][22]  ( .D(
        write_data_reg[22]), .E(n6844), .C(n1107), .RN(n6621), .Q(n5834) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][24]  ( .D(
        write_data_reg[24]), .E(n6844), .C(n1107), .RN(n6621), .Q(n5861) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][25]  ( .D(n6981), .E(
        n6843), .C(n1107), .RN(n6621), .Q(n5915) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][26]  ( .D(n6983), .E(
        n6843), .C(n1107), .RN(n6621), .Q(n5909) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][27]  ( .D(n6985), .E(
        n6843), .C(n1107), .RN(n6621), .Q(n5914) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][28]  ( .D(n6987), .E(
        n6843), .C(n1107), .RN(n6621), .Q(n5912) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][29]  ( .D(n6989), .E(
        n6843), .C(n1107), .RN(n6621), .Q(n5911) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][30]  ( .D(n6991), .E(
        n6843), .C(n1107), .RN(n6622), .Q(n5913) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[16][31]  ( .D(n6993), .E(
        n6843), .C(n1107), .RN(n6622), .Q(n6021) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][0]  ( .D(
        write_data_reg[0]), .E(n6857), .C(n1107), .RN(n6638), .Q(n6039) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][1]  ( .D(n6932), .E(
        n6857), .C(n1107), .RN(n6638), .Q(n6038) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][2]  ( .D(n6934), .E(
        n6857), .C(n1107), .RN(n6638), .Q(n6023) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][3]  ( .D(n6937), .E(
        n6857), .C(n1107), .RN(n6638), .Q(n6037) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][4]  ( .D(
        write_data_reg[4]), .E(n6856), .C(n1107), .RN(n6639), .Q(n6036) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][5]  ( .D(
        write_data_reg[5]), .E(n6856), .C(n1107), .RN(n6639), .Q(n5927) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][6]  ( .D(
        write_data_reg[6]), .E(n6856), .C(n1107), .RN(n6639), .Q(n5842) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][9]  ( .D(n6949), .E(
        n6856), .C(n1107), .RN(n6639), .Q(n6041) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][10]  ( .D(n6951), .E(
        n6856), .C(n1107), .RN(n6639), .Q(n6035) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][17]  ( .D(n6965), .E(
        n6855), .C(n1107), .RN(n6640), .Q(n6032) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][18]  ( .D(n6967), .E(
        n6854), .C(n1107), .RN(n6640), .Q(n5940) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][20]  ( .D(n6971), .E(
        n6854), .C(n1107), .RN(n6640), .Q(n5916) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][21]  ( .D(n6973), .E(
        n6854), .C(n1107), .RN(n6640), .Q(n5864) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][22]  ( .D(
        write_data_reg[22]), .E(n6854), .C(n1107), .RN(n6641), .Q(n5836) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][23]  ( .D(n6977), .E(
        n6854), .C(n1107), .RN(n6641), .Q(n6040) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][24]  ( .D(
        write_data_reg[24]), .E(n6854), .C(n1107), .RN(n6641), .Q(n5862) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][25]  ( .D(n6981), .E(
        n6853), .C(n1107), .RN(n6641), .Q(n6028) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][26]  ( .D(n6983), .E(
        n6853), .C(n1107), .RN(n6641), .Q(n5908) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][27]  ( .D(n6985), .E(
        n6853), .C(n1107), .RN(n6641), .Q(n6027) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][28]  ( .D(n6987), .E(
        n6853), .C(n1107), .RN(n6641), .Q(n6025) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][29]  ( .D(n6989), .E(
        n6853), .C(n1107), .RN(n6641), .Q(n6024) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][30]  ( .D(n6991), .E(
        n6853), .C(n1107), .RN(n6641), .Q(n6026) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[18][31]  ( .D(n6993), .E(
        n6853), .C(n1107), .RN(n6642), .Q(n6022) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][1]  ( .D(
        write_data_reg[1]), .E(n6862), .C(n1107), .RN(n6666), .Q(n6059) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][2]  ( .D(
        write_data_reg[2]), .E(n6862), .C(n1107), .RN(n6666), .Q(n6043) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][25]  ( .D(n6981), .E(
        n6858), .C(n1107), .RN(n6669), .Q(n6048) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][26]  ( .D(n6983), .E(
        n6858), .C(n1107), .RN(n6669), .Q(n6042) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][27]  ( .D(n6985), .E(
        n6858), .C(n1107), .RN(n6669), .Q(n6047) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][28]  ( .D(n6987), .E(
        n6858), .C(n1107), .RN(n6669), .Q(n6045) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][29]  ( .D(n6989), .E(
        n6858), .C(n1107), .RN(n6669), .Q(n6044) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][30]  ( .D(n6991), .E(
        n6858), .C(n1107), .RN(n6669), .Q(n6046) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[19][31]  ( .D(
        write_data_reg[31]), .E(n6858), .C(n1107), .RN(n6669), .Q(n5932) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][1]  ( .D(
        write_data_reg[1]), .E(n6882), .C(n1107), .RN(n6694), .QN(n6006) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][2]  ( .D(
        write_data_reg[2]), .E(n6882), .C(n1107), .RN(n6694), .QN(n6066) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][6]  ( .D(n6943), .E(
        n6881), .C(n1107), .RN(n6695), .QN(n6014) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][22]  ( .D(n6975), .E(
        n6879), .C(n1107), .RN(n6696), .QN(n6008) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][24]  ( .D(n6979), .E(
        n6879), .C(n1107), .RN(n6696), .QN(n6009) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][25]  ( .D(n6981), .E(
        n6879), .C(n1107), .RN(n6697), .QN(n5903) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][26]  ( .D(
        write_data_reg[26]), .E(n6879), .C(n1107), .RN(n6697), .QN(n6063) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][29]  ( .D(n6989), .E(
        n6878), .C(n1107), .RN(n6697), .QN(n6065) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][30]  ( .D(n6991), .E(
        n6878), .C(n1107), .RN(n6697), .QN(n6062) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][31]  ( .D(
        write_data_reg[31]), .E(n6878), .C(n1107), .RN(n6697), .QN(n5939) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][0]  ( .D(
        write_data_reg[0]), .E(n6872), .C(n1107), .RN(n6697), .QN(n5974) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][1]  ( .D(n6932), .E(
        n6872), .C(n1107), .RN(n6697), .QN(n5981) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][2]  ( .D(n6934), .E(
        n6872), .C(n1107), .RN(n6697), .QN(n5989) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][3]  ( .D(n6936), .E(
        n6872), .C(n1107), .RN(n6697), .QN(n5991) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][4]  ( .D(n6939), .E(
        n6871), .C(n1107), .RN(n6698), .QN(n5992) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][5]  ( .D(n6941), .E(
        n6871), .C(n1107), .RN(n6698), .QN(n5993) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][6]  ( .D(n6943), .E(
        n6871), .C(n1107), .RN(n6698), .QN(n5994) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][8]  ( .D(n6947), .E(
        n6871), .C(n1107), .RN(n6698), .QN(n5996) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][9]  ( .D(n6949), .E(
        n6871), .C(n1107), .RN(n6698), .QN(n5997) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][10]  ( .D(
        write_data_reg[10]), .E(n6871), .C(n1107), .RN(n6698), .QN(n5975) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][14]  ( .D(
        write_data_reg[14]), .E(n6870), .C(n1107), .RN(n6699), .QN(n5978) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][16]  ( .D(n6963), .E(
        n6870), .C(n1107), .RN(n6699), .QN(n5980) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][17]  ( .D(
        write_data_reg[17]), .E(n6870), .C(n1107), .RN(n6699), .QN(n5882) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][18]  ( .D(n6967), .E(
        n6869), .C(n1107), .RN(n6699), .QN(n5874) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][19]  ( .D(
        write_data_reg[19]), .E(n6869), .C(n1107), .RN(n6699), .QN(n5883) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][20]  ( .D(
        write_data_reg[20]), .E(n6869), .C(n1107), .RN(n6699), .QN(n5884) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][21]  ( .D(
        write_data_reg[21]), .E(n6869), .C(n1107), .RN(n6699), .QN(n5982) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][22]  ( .D(n6975), .E(
        n6869), .C(n1107), .RN(n6700), .QN(n5983) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][23]  ( .D(
        write_data_reg[23]), .E(n6869), .C(n1107), .RN(n6700), .QN(n5886) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][24]  ( .D(n6979), .E(
        n6869), .C(n1107), .RN(n6700), .QN(n5887) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][25]  ( .D(n6981), .E(
        n6868), .C(n1107), .RN(n6700), .QN(n5984) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][26]  ( .D(
        write_data_reg[26]), .E(n6868), .C(n1107), .RN(n6700), .QN(n5985) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][28]  ( .D(n6987), .E(
        n6868), .C(n1107), .RN(n6700), .QN(n5987) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][29]  ( .D(n6989), .E(
        n6868), .C(n1107), .RN(n6700), .QN(n5988) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][30]  ( .D(n6991), .E(
        n6868), .C(n1107), .RN(n6700), .QN(n5990) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][31]  ( .D(
        write_data_reg[31]), .E(n6868), .C(n1107), .RN(n6700), .QN(n5890) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][0]  ( .D(
        write_data_reg[0]), .E(n6792), .C(n1107), .RN(n6706), .QN(n5947) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][1]  ( .D(
        write_data_reg[1]), .E(n6792), .C(n1107), .RN(n6706), .QN(n5954) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][2]  ( .D(
        write_data_reg[2]), .E(n6792), .C(n1107), .RN(n6707), .QN(n5963) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][3]  ( .D(n6936), .E(n6792), .C(n1107), .RN(n6707), .QN(n5965) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][4]  ( .D(
        write_data_reg[4]), .E(n6791), .C(n1107), .RN(n6707), .QN(n5966) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][5]  ( .D(n6941), .E(n6791), .C(n1107), .RN(n6707), .QN(n5967) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][6]  ( .D(n6943), .E(n6791), .C(n1107), .RN(n6707), .QN(n5968) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][7]  ( .D(n6945), .E(n6791), .C(n1107), .RN(n6707), .QN(n5969) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][8]  ( .D(n6947), .E(n6791), .C(n1107), .RN(n6707), .QN(n5970) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][9]  ( .D(n6949), .E(n6791), .C(n1107), .RN(n6707), .QN(n5971) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][10]  ( .D(
        write_data_reg[10]), .E(n6791), .C(n1107), .RN(n6707), .QN(n5948) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][12]  ( .D(
        write_data_reg[12]), .E(n6790), .C(n1107), .RN(n6708), .QN(n5950) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][13]  ( .D(n6957), .E(
        n6790), .C(n1107), .RN(n6708), .QN(n5972) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][14]  ( .D(
        write_data_reg[14]), .E(n6790), .C(n1107), .RN(n6708), .QN(n5951) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][15]  ( .D(n6961), .E(
        n6790), .C(n1107), .RN(n6708), .QN(n5952) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][16]  ( .D(n6963), .E(
        n6790), .C(n1107), .RN(n6708), .QN(n5953) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][17]  ( .D(
        write_data_reg[17]), .E(n6790), .C(n1107), .RN(n6708), .QN(n5869) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][18]  ( .D(n6967), .E(
        n6790), .C(n1107), .RN(n6708), .QN(n5973) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][20]  ( .D(
        write_data_reg[20]), .E(n6789), .C(n1107), .RN(n6708), .QN(n5871) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][21]  ( .D(
        write_data_reg[21]), .E(n6789), .C(n1107), .RN(n6708), .QN(n5955) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][22]  ( .D(n6975), .E(
        n6789), .C(n1107), .RN(n6709), .QN(n5956) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][24]  ( .D(n6979), .E(
        n6789), .C(n1107), .RN(n6709), .QN(n5957) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][25]  ( .D(n6981), .E(
        n6789), .C(n1107), .RN(n6709), .QN(n5958) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][26]  ( .D(
        write_data_reg[26]), .E(n6789), .C(n1107), .RN(n6709), .QN(n5959) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][29]  ( .D(n6989), .E(
        n6789), .C(n1107), .RN(n6709), .QN(n5962) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][30]  ( .D(n6991), .E(
        n6788), .C(n1107), .RN(n6709), .QN(n5964) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][31]  ( .D(
        write_data_reg[31]), .E(n6788), .C(n1107), .RN(n6709), .QN(n5873) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][1]  ( .D(n6932), .E(
        n6877), .C(n1107), .RN(n6713), .QN(n5839) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][2]  ( .D(n6934), .E(
        n6877), .C(n1107), .RN(n6713), .QN(n5840) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][4]  ( .D(n6939), .E(
        n6876), .C(n1107), .RN(n6713), .QN(n5892) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][5]  ( .D(n6941), .E(
        n6876), .C(n1107), .RN(n6713), .QN(n5893) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][6]  ( .D(n6943), .E(
        n6876), .C(n1107), .RN(n6713), .QN(n5894) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][9]  ( .D(n6949), .E(
        n6876), .C(n1107), .RN(n6714), .QN(n5857) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][10]  ( .D(
        write_data_reg[10]), .E(n6876), .C(n1107), .RN(n6714), .QN(n5876) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][18]  ( .D(n6967), .E(
        n6874), .C(n1107), .RN(n6715), .QN(n5875) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][20]  ( .D(
        write_data_reg[20]), .E(n6874), .C(n1107), .RN(n6715), .QN(n5853) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][21]  ( .D(
        write_data_reg[21]), .E(n6874), .C(n1107), .RN(n6715), .QN(n5885) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][22]  ( .D(n6975), .E(
        n6874), .C(n1107), .RN(n6715), .QN(n5854) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][23]  ( .D(
        write_data_reg[23]), .E(n6874), .C(n1107), .RN(n6715), .QN(n5855) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][24]  ( .D(n6979), .E(
        n6874), .C(n1107), .RN(n6715), .QN(n5888) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][25]  ( .D(n6981), .E(
        n6873), .C(n1107), .RN(n6716), .QN(n5856) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][26]  ( .D(
        write_data_reg[26]), .E(n6873), .C(n1107), .RN(n6716), .QN(n5905) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][27]  ( .D(n6985), .E(
        n6873), .C(n1107), .RN(n6716), .QN(n5889) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][28]  ( .D(n6987), .E(
        n6873), .C(n1107), .RN(n6716), .QN(n5906) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][29]  ( .D(n6989), .E(
        n6873), .C(n1107), .RN(n6716), .QN(n5907) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][30]  ( .D(n6991), .E(
        n6873), .C(n1107), .RN(n6716), .QN(n5904) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][31]  ( .D(
        write_data_reg[31]), .E(n6873), .C(n1107), .RN(n6716), .QN(n5858) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][27]  ( .D(n6985), .E(
        n6878), .C(n1107), .RN(n6720), .QN(n6010) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[23][28]  ( .D(n6987), .E(
        n6878), .C(n1107), .RN(n6720), .QN(n6064) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[21][27]  ( .D(n6985), .E(
        n6868), .C(n1107), .RN(n6721), .QN(n5986) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][19]  ( .D(
        write_data_reg[19]), .E(n6788), .C(n1107), .RN(n6722), .QN(n5870) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][23]  ( .D(
        write_data_reg[23]), .E(n6788), .C(n1107), .RN(n6722), .QN(n5872) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][27]  ( .D(n6985), .E(
        n6788), .C(n1107), .RN(n6722), .QN(n5960) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[5][28]  ( .D(n6987), .E(
        n6788), .C(n1107), .RN(n6722), .QN(n5961) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][14]  ( .D(
        write_data_reg[14]), .E(n6823), .C(n1107), .RN(n6725), .QN(n5081) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][8]  ( .D(n6947), .E(
        n6833), .C(n1107), .RN(n6724), .QN(n4939) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][18]  ( .D(n6967), .E(
        n6833), .C(n1107), .RN(n6724), .QN(n4891) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][4]  ( .D(n6939), .E(
        n6834), .C(n1107), .RN(n6724), .QN(n4945) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][26]  ( .D(
        write_data_reg[26]), .E(n6833), .C(n1107), .RN(n6723), .QN(n4877) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][23]  ( .D(
        write_data_reg[23]), .E(n6888), .C(n1107), .RN(n6723), .QN(n4883) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][24]  ( .D(n6979), .E(
        n6833), .C(n1107), .RN(n6723), .QN(n5325) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][27]  ( .D(n6985), .E(
        n6898), .C(n1107), .RN(n6724), .QN(n5021) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][27]  ( .D(n6985), .E(
        n6833), .C(n1107), .RN(n6723), .QN(n4915) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][13]  ( .D(n6957), .E(
        n6834), .C(n1107), .RN(n6724), .QN(n4907) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][4]  ( .D(n6939), .E(n6898), .C(n1107), .RN(n6724), .QN(n5327) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][23]  ( .D(
        write_data_reg[23]), .E(n6833), .C(n1107), .RN(n6724), .QN(n4931) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][10]  ( .D(
        write_data_reg[10]), .E(n6834), .C(n1107), .RN(n6724), .QN(n4905) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][14]  ( .D(
        write_data_reg[14]), .E(n6833), .C(n1107), .RN(n6724), .QN(n4885) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][22]  ( .D(
        write_data_reg[22]), .E(n6902), .C(n1107), .RN(n6611), .QN(n5337) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][0]  ( .D(
        write_data_reg[0]), .E(n6827), .C(n1107), .RN(n6611), .QN(n5287) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][1]  ( .D(
        write_data_reg[1]), .E(n6827), .C(n1107), .RN(n6611), .QN(n5299) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][2]  ( .D(
        write_data_reg[2]), .E(n6827), .C(n1107), .RN(n6611), .QN(n5195) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][3]  ( .D(n6937), .E(
        n6827), .C(n1107), .RN(n6612), .QN(n5281) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][4]  ( .D(
        write_data_reg[4]), .E(n6826), .C(n1107), .RN(n6612), .QN(n5271) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][5]  ( .D(
        write_data_reg[5]), .E(n6826), .C(n1107), .RN(n6612), .QN(n5235) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][6]  ( .D(
        write_data_reg[6]), .E(n6826), .C(n1107), .RN(n6612), .QN(n5189) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][7]  ( .D(
        write_data_reg[7]), .E(n6826), .C(n1107), .RN(n6612), .QN(n5275) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][8]  ( .D(n6947), .E(
        n6826), .C(n1107), .RN(n6612), .QN(n5253) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][9]  ( .D(n6949), .E(
        n6826), .C(n1107), .RN(n6612), .QN(n5201) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][10]  ( .D(
        write_data_reg[10]), .E(n6826), .C(n1107), .RN(n6612), .QN(n5145) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][11]  ( .D(
        write_data_reg[11]), .E(n6825), .C(n1107), .RN(n6612), .QN(n5247) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][12]  ( .D(n6955), .E(
        n6825), .C(n1107), .RN(n6613), .QN(n5207) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][13]  ( .D(n6957), .E(
        n6825), .C(n1107), .RN(n6613), .QN(n5151) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][15]  ( .D(
        write_data_reg[15]), .E(n6825), .C(n1107), .RN(n6613), .QN(n5265) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][16]  ( .D(
        write_data_reg[16]), .E(n6825), .C(n1107), .RN(n6613), .QN(n5223) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][17]  ( .D(n6965), .E(
        n6825), .C(n1107), .RN(n6613), .QN(n5167) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][18]  ( .D(n6967), .E(
        n6825), .C(n1107), .RN(n6613), .QN(n5105) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][19]  ( .D(n6969), .E(
        n6824), .C(n1107), .RN(n6613), .QN(n5259) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][20]  ( .D(n6971), .E(
        n6824), .C(n1107), .RN(n6613), .QN(n5217) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][21]  ( .D(n6973), .E(
        n6824), .C(n1107), .RN(n6613), .QN(n5161) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][22]  ( .D(
        write_data_reg[22]), .E(n6824), .C(n1107), .RN(n6614), .QN(n5093) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][23]  ( .D(
        write_data_reg[23]), .E(n6824), .C(n1107), .RN(n6614), .QN(n5229) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][24]  ( .D(n6979), .E(
        n6824), .C(n1107), .RN(n6614), .QN(n5183) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][25]  ( .D(n6981), .E(
        n6824), .C(n1107), .RN(n6614), .QN(n5129) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][26]  ( .D(
        write_data_reg[26]), .E(n6823), .C(n1107), .RN(n6614), .QN(n5057) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][27]  ( .D(n6985), .E(
        n6823), .C(n1107), .RN(n6614), .QN(n5173) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][28]  ( .D(n6987), .E(
        n6823), .C(n1107), .RN(n6614), .QN(n5117) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][29]  ( .D(n6989), .E(
        n6823), .C(n1107), .RN(n6614), .QN(n5041) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][30]  ( .D(n6991), .E(
        n6823), .C(n1107), .RN(n6614), .QN(n4991) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[28][31]  ( .D(n6993), .E(
        n6823), .C(n1107), .RN(n6615), .QN(n5241) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][0]  ( .D(n6930), .E(
        n6807), .C(n1107), .RN(n6615), .QN(n5291) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][1]  ( .D(
        write_data_reg[1]), .E(n6807), .C(n1107), .RN(n6615), .QN(n5303) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][2]  ( .D(
        write_data_reg[2]), .E(n6807), .C(n1107), .RN(n6615), .QN(n5199) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][3]  ( .D(n6937), .E(
        n6807), .C(n1107), .RN(n6615), .QN(n5285) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][4]  ( .D(
        write_data_reg[4]), .E(n6806), .C(n1107), .RN(n6615), .QN(n5345) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][5]  ( .D(
        write_data_reg[5]), .E(n6806), .C(n1107), .RN(n6615), .QN(n5239) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][6]  ( .D(
        write_data_reg[6]), .E(n6806), .C(n1107), .RN(n6615), .QN(n5193) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][7]  ( .D(
        write_data_reg[7]), .E(n6806), .C(n1107), .RN(n6615), .QN(n5279) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][8]  ( .D(
        write_data_reg[8]), .E(n6806), .C(n1107), .RN(n6616), .QN(n5257) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][9]  ( .D(n6949), .E(
        n6806), .C(n1107), .RN(n6616), .QN(n5205) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][10]  ( .D(n6951), .E(
        n6806), .C(n1107), .RN(n6616), .QN(n5149) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][11]  ( .D(
        write_data_reg[11]), .E(n6805), .C(n1107), .RN(n6616), .QN(n5251) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][12]  ( .D(n6955), .E(
        n6805), .C(n1107), .RN(n6616), .QN(n5211) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][13]  ( .D(
        write_data_reg[13]), .E(n6805), .C(n1107), .RN(n6616), .QN(n5155) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][14]  ( .D(
        write_data_reg[14]), .E(n6805), .C(n1107), .RN(n6616), .QN(n5085) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][15]  ( .D(
        write_data_reg[15]), .E(n6805), .C(n1107), .RN(n6616), .QN(n5269) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][16]  ( .D(
        write_data_reg[16]), .E(n6805), .C(n1107), .RN(n6616), .QN(n5227) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][17]  ( .D(n6965), .E(
        n6805), .C(n1107), .RN(n6617), .QN(n5171) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][18]  ( .D(n6967), .E(
        n6804), .C(n1107), .RN(n6617), .QN(n5109) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][19]  ( .D(n6969), .E(
        n6804), .C(n1107), .RN(n6617), .QN(n5263) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][20]  ( .D(n6971), .E(
        n6804), .C(n1107), .RN(n6617), .QN(n5221) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][21]  ( .D(n6973), .E(
        n6804), .C(n1107), .RN(n6617), .QN(n5165) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][22]  ( .D(
        write_data_reg[22]), .E(n6804), .C(n1107), .RN(n6617), .QN(n5097) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][23]  ( .D(n6977), .E(
        n6804), .C(n1107), .RN(n6617), .QN(n5233) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][24]  ( .D(
        write_data_reg[24]), .E(n6804), .C(n1107), .RN(n6617), .QN(n5187) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][25]  ( .D(n6981), .E(
        n6803), .C(n1107), .RN(n6617), .QN(n5343) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][26]  ( .D(n6983), .E(
        n6803), .C(n1107), .RN(n6618), .QN(n5061) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][27]  ( .D(n6985), .E(
        n6803), .C(n1107), .RN(n6618), .QN(n5335) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][28]  ( .D(n6987), .E(
        n6803), .C(n1107), .RN(n6618), .QN(n5121) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][29]  ( .D(n6989), .E(
        n6803), .C(n1107), .RN(n6618), .QN(n5045) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][31]  ( .D(n6993), .E(
        n6803), .C(n1107), .RN(n6618), .QN(n5245) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][0]  ( .D(
        write_data_reg[0]), .E(n6922), .C(n1107), .RN(n6622), .QN(n4949) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][1]  ( .D(
        write_data_reg[1]), .E(n6922), .C(n1107), .RN(n6622), .QN(n5293) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][2]  ( .D(
        write_data_reg[2]), .E(n6922), .C(n1107), .RN(n6622), .QN(n5035) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][3]  ( .D(n6937), .E(
        n6922), .C(n1107), .RN(n6622), .QN(n5213) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][4]  ( .D(
        write_data_reg[4]), .E(n6921), .C(n1107), .RN(n6622), .QN(n5157) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][5]  ( .D(
        write_data_reg[5]), .E(n6921), .C(n1107), .RN(n6622), .QN(n5087) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][6]  ( .D(
        write_data_reg[6]), .E(n6921), .C(n1107), .RN(n6622), .QN(n5029) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][7]  ( .D(
        write_data_reg[7]), .E(n6921), .C(n1107), .RN(n6623), .QN(n5177) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][8]  ( .D(
        write_data_reg[8]), .E(n6921), .C(n1107), .RN(n6623), .QN(n5123) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][9]  ( .D(n6949), .E(
        n6921), .C(n1107), .RN(n6623), .QN(n5047) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][10]  ( .D(n6951), .E(
        n6921), .C(n1107), .RN(n6623), .QN(n4997) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][11]  ( .D(
        write_data_reg[11]), .E(n6920), .C(n1107), .RN(n6623), .QN(n5111) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][12]  ( .D(n6955), .E(
        n6920), .C(n1107), .RN(n6623), .QN(n5051) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][13]  ( .D(
        write_data_reg[13]), .E(n6920), .C(n1107), .RN(n6623), .QN(n5001) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][14]  ( .D(n6959), .E(
        n6920), .C(n1107), .RN(n6623), .QN(n4969) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][15]  ( .D(
        write_data_reg[15]), .E(n6920), .C(n1107), .RN(n6623), .QN(n5139) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][16]  ( .D(
        write_data_reg[16]), .E(n6920), .C(n1107), .RN(n6624), .QN(n5069) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][17]  ( .D(n6965), .E(
        n6920), .C(n1107), .RN(n6624), .QN(n5011) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][18]  ( .D(n6967), .E(
        n6919), .C(n1107), .RN(n6624), .QN(n4977) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][19]  ( .D(n6969), .E(
        n6919), .C(n1107), .RN(n6624), .QN(n5133) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][20]  ( .D(n6971), .E(
        n6919), .C(n1107), .RN(n6624), .QN(n5063) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][21]  ( .D(n6973), .E(
        n6919), .C(n1107), .RN(n6624), .QN(n5007) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][22]  ( .D(
        write_data_reg[22]), .E(n6919), .C(n1107), .RN(n6624), .QN(n4973) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][23]  ( .D(n6977), .E(
        n6919), .C(n1107), .RN(n6624), .QN(n5075) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][24]  ( .D(
        write_data_reg[24]), .E(n6919), .C(n1107), .RN(n6624), .QN(n5023) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][25]  ( .D(n6981), .E(
        n6918), .C(n1107), .RN(n6625), .QN(n4987) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][26]  ( .D(n6983), .E(
        n6918), .C(n1107), .RN(n6625), .QN(n4965) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][27]  ( .D(n6985), .E(
        n6918), .C(n1107), .RN(n6625), .QN(n5017) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][28]  ( .D(n6987), .E(
        n6918), .C(n1107), .RN(n6625), .QN(n4983) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][29]  ( .D(n6989), .E(
        n6918), .C(n1107), .RN(n6625), .QN(n4959) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][30]  ( .D(n6991), .E(
        n6918), .C(n1107), .RN(n6625), .QN(n4953) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[12][31]  ( .D(n6993), .E(
        n6918), .C(n1107), .RN(n6625), .QN(n5099) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][0]  ( .D(n6930), .E(n6902), .C(n1107), .RN(n6625), .QN(n5315) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][1]  ( .D(
        write_data_reg[1]), .E(n6902), .C(n1107), .RN(n6625), .QN(n5297) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][2]  ( .D(
        write_data_reg[2]), .E(n6902), .C(n1107), .RN(n6626), .QN(n5039) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][3]  ( .D(n6937), .E(n6901), .C(n1107), .RN(n6626), .QN(n5317) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][5]  ( .D(
        write_data_reg[5]), .E(n6901), .C(n1107), .RN(n6626), .QN(n5091) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][6]  ( .D(
        write_data_reg[6]), .E(n6901), .C(n1107), .RN(n6626), .QN(n5033) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][7]  ( .D(
        write_data_reg[7]), .E(n6901), .C(n1107), .RN(n6626), .QN(n5181) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][8]  ( .D(
        write_data_reg[8]), .E(n6901), .C(n1107), .RN(n6626), .QN(n5127) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][9]  ( .D(n6949), .E(n6901), .C(n1107), .RN(n6626), .QN(n5341) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][10]  ( .D(n6951), .E(
        n6901), .C(n1107), .RN(n6626), .QN(n5349) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][11]  ( .D(
        write_data_reg[11]), .E(n6900), .C(n1107), .RN(n6626), .QN(n5115) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][12]  ( .D(n6955), .E(
        n6900), .C(n1107), .RN(n6627), .QN(n5055) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][13]  ( .D(
        write_data_reg[13]), .E(n6900), .C(n1107), .RN(n6627), .QN(n5005) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][14]  ( .D(n6959), .E(
        n6900), .C(n1107), .RN(n6627), .QN(n5313) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][15]  ( .D(
        write_data_reg[15]), .E(n6900), .C(n1107), .RN(n6627), .QN(n5143) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][16]  ( .D(
        write_data_reg[16]), .E(n6900), .C(n1107), .RN(n6627), .QN(n5073) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][17]  ( .D(n6965), .E(
        n6900), .C(n1107), .RN(n6627), .QN(n5015) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][18]  ( .D(n6967), .E(
        n6899), .C(n1107), .RN(n6627), .QN(n4981) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][19]  ( .D(n6969), .E(
        n6899), .C(n1107), .RN(n6627), .QN(n5137) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][20]  ( .D(n6971), .E(
        n6899), .C(n1107), .RN(n6627), .QN(n5067) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][21]  ( .D(n6973), .E(
        n6899), .C(n1107), .RN(n6628), .QN(n5323) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][23]  ( .D(n6977), .E(
        n6899), .C(n1107), .RN(n6628), .QN(n5079) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][24]  ( .D(
        write_data_reg[24]), .E(n6899), .C(n1107), .RN(n6628), .QN(n5027) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][25]  ( .D(n6981), .E(
        n6899), .C(n1107), .RN(n6628), .QN(n5333) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][26]  ( .D(n6983), .E(
        n6898), .C(n1107), .RN(n6628), .QN(n5339) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][28]  ( .D(n6987), .E(
        n6898), .C(n1107), .RN(n6628), .QN(n5351) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][29]  ( .D(n6989), .E(
        n6898), .C(n1107), .RN(n6628), .QN(n4963) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][30]  ( .D(n6991), .E(
        n6898), .C(n1107), .RN(n6628), .QN(n4957) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[8][31]  ( .D(n6993), .E(
        n6898), .C(n1107), .RN(n6628), .QN(n5103) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][0]  ( .D(
        write_data_reg[0]), .E(n6767), .C(n1107), .RN(n6629), .QN(n4707) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][1]  ( .D(
        write_data_reg[1]), .E(n6767), .C(n1107), .RN(n6629), .QN(n4663) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][2]  ( .D(
        write_data_reg[2]), .E(n6767), .C(n1107), .RN(n6629), .QN(n4659) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][3]  ( .D(n6937), .E(n6767), .C(n1107), .RN(n6629), .QN(n4655) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][4]  ( .D(
        write_data_reg[4]), .E(n6766), .C(n1107), .RN(n6629), .QN(n4651) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][5]  ( .D(
        write_data_reg[5]), .E(n6766), .C(n1107), .RN(n6629), .QN(n4647) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][6]  ( .D(
        write_data_reg[6]), .E(n6766), .C(n1107), .RN(n6629), .QN(n4643) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][7]  ( .D(
        write_data_reg[7]), .E(n6766), .C(n1107), .RN(n6629), .QN(n4639) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][8]  ( .D(
        write_data_reg[8]), .E(n6766), .C(n1107), .RN(n6629), .QN(n4635) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][9]  ( .D(n6949), .E(n6766), .C(n1107), .RN(n6630), .QN(n4631) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][10]  ( .D(n6951), .E(
        n6766), .C(n1107), .RN(n6630), .QN(n4703) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][11]  ( .D(
        write_data_reg[11]), .E(n6765), .C(n1107), .RN(n6630), .QN(n4699) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][12]  ( .D(n6955), .E(
        n6765), .C(n1107), .RN(n6630), .QN(n4695) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][13]  ( .D(
        write_data_reg[13]), .E(n6765), .C(n1107), .RN(n6630), .QN(n4691) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][14]  ( .D(n6959), .E(
        n6765), .C(n1107), .RN(n6630), .QN(n4687) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][15]  ( .D(
        write_data_reg[15]), .E(n6765), .C(n1107), .RN(n6630), .QN(n4683) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][16]  ( .D(
        write_data_reg[16]), .E(n6765), .C(n1107), .RN(n6630), .QN(n4679) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][17]  ( .D(n6965), .E(
        n6765), .C(n1107), .RN(n6630), .QN(n4675) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][18]  ( .D(n6967), .E(
        n6764), .C(n1107), .RN(n6631), .QN(n4671) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][19]  ( .D(n6969), .E(
        n6764), .C(n1107), .RN(n6631), .QN(n4667) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][20]  ( .D(n6971), .E(
        n6764), .C(n1107), .RN(n6631), .QN(n4627) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][21]  ( .D(n6973), .E(
        n6764), .C(n1107), .RN(n6631), .QN(n4623) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][22]  ( .D(
        write_data_reg[22]), .E(n6764), .C(n1107), .RN(n6631), .QN(n4619) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][23]  ( .D(n6977), .E(
        n6764), .C(n1107), .RN(n6631), .QN(n4615) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][24]  ( .D(
        write_data_reg[24]), .E(n6764), .C(n1107), .RN(n6631), .QN(n4611) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][25]  ( .D(n6981), .E(
        n6763), .C(n1107), .RN(n6631), .QN(n4607) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][26]  ( .D(n6983), .E(
        n6763), .C(n1107), .RN(n6631), .QN(n4603) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][27]  ( .D(n6985), .E(
        n6763), .C(n1107), .RN(n6632), .QN(n4599) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][28]  ( .D(n6987), .E(
        n6763), .C(n1107), .RN(n6632), .QN(n4595) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][29]  ( .D(n6989), .E(
        n6763), .C(n1107), .RN(n6632), .QN(n4591) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][30]  ( .D(n6991), .E(
        n6763), .C(n1107), .RN(n6632), .QN(n4587) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[0][31]  ( .D(n6993), .E(
        n6763), .C(n1107), .RN(n6632), .QN(n4583) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][0]  ( .D(n6930), .E(
        n6837), .C(n1107), .RN(n6632), .QN(n5331) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][1]  ( .D(
        write_data_reg[1]), .E(n6837), .C(n1107), .RN(n6632), .QN(n5305) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][2]  ( .D(
        write_data_reg[2]), .E(n6837), .C(n1107), .RN(n6632), .QN(n4921) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][3]  ( .D(n6937), .E(
        n6837), .C(n1107), .RN(n6632), .QN(n5321) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][5]  ( .D(
        write_data_reg[5]), .E(n6836), .C(n1107), .RN(n6633), .QN(n4933) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][6]  ( .D(
        write_data_reg[6]), .E(n6836), .C(n1107), .RN(n6633), .QN(n4919) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][7]  ( .D(
        write_data_reg[7]), .E(n6836), .C(n1107), .RN(n6633), .QN(n4947) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][9]  ( .D(n6949), .E(
        n6836), .C(n1107), .RN(n6633), .QN(n5319) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][11]  ( .D(
        write_data_reg[11]), .E(n6836), .C(n1107), .RN(n6633), .QN(n4937) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][12]  ( .D(n6955), .E(
        n6836), .C(n1107), .RN(n6633), .QN(n4923) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][15]  ( .D(
        write_data_reg[15]), .E(n6836), .C(n1107), .RN(n6633), .QN(n4943) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][16]  ( .D(
        write_data_reg[16]), .E(n6835), .C(n1107), .RN(n6633), .QN(n4929) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][17]  ( .D(n6965), .E(
        n6835), .C(n1107), .RN(n6633), .QN(n4913) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][19]  ( .D(n6969), .E(
        n6835), .C(n1107), .RN(n6634), .QN(n4941) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][20]  ( .D(n6971), .E(
        n6835), .C(n1107), .RN(n6634), .QN(n4927) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][21]  ( .D(n6973), .E(
        n6835), .C(n1107), .RN(n6634), .QN(n4911) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][22]  ( .D(
        write_data_reg[22]), .E(n6835), .C(n1107), .RN(n6634), .QN(n5329) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][25]  ( .D(n6981), .E(
        n6835), .C(n1107), .RN(n6634), .QN(n4899) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][28]  ( .D(n6987), .E(
        n6834), .C(n1107), .RN(n6634), .QN(n4895) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][29]  ( .D(n6989), .E(
        n6834), .C(n1107), .RN(n6634), .QN(n4871) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][30]  ( .D(n6991), .E(
        n6834), .C(n1107), .RN(n6634), .QN(n4853) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[30][31]  ( .D(n6993), .E(
        n6834), .C(n1107), .RN(n6634), .QN(n4935) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][0]  ( .D(
        write_data_reg[0]), .E(n6817), .C(n1107), .RN(n6635), .QN(n5289) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][1]  ( .D(
        write_data_reg[1]), .E(n6817), .C(n1107), .RN(n6635), .QN(n5301) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][2]  ( .D(
        write_data_reg[2]), .E(n6817), .C(n1107), .RN(n6635), .QN(n5197) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][3]  ( .D(n6937), .E(
        n6817), .C(n1107), .RN(n6635), .QN(n5283) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][4]  ( .D(
        write_data_reg[4]), .E(n6816), .C(n1107), .RN(n6635), .QN(n5273) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][5]  ( .D(
        write_data_reg[5]), .E(n6816), .C(n1107), .RN(n6635), .QN(n5237) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][6]  ( .D(
        write_data_reg[6]), .E(n6816), .C(n1107), .RN(n6635), .QN(n5191) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][7]  ( .D(
        write_data_reg[7]), .E(n6816), .C(n1107), .RN(n6635), .QN(n5277) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][8]  ( .D(
        write_data_reg[8]), .E(n6816), .C(n1107), .RN(n6635), .QN(n5255) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][9]  ( .D(n6949), .E(
        n6816), .C(n1107), .RN(n6636), .QN(n5203) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][10]  ( .D(n6951), .E(
        n6816), .C(n1107), .RN(n6636), .QN(n5147) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][11]  ( .D(
        write_data_reg[11]), .E(n6815), .C(n1107), .RN(n6636), .QN(n5249) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][12]  ( .D(n6955), .E(
        n6815), .C(n1107), .RN(n6636), .QN(n5209) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][13]  ( .D(
        write_data_reg[13]), .E(n6815), .C(n1107), .RN(n6636), .QN(n5153) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][14]  ( .D(n6959), .E(
        n6815), .C(n1107), .RN(n6636), .QN(n5083) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][15]  ( .D(
        write_data_reg[15]), .E(n6815), .C(n1107), .RN(n6636), .QN(n5267) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][16]  ( .D(
        write_data_reg[16]), .E(n6815), .C(n1107), .RN(n6636), .QN(n5225) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][17]  ( .D(n6965), .E(
        n6815), .C(n1107), .RN(n6636), .QN(n5169) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][18]  ( .D(n6967), .E(
        n6814), .C(n1107), .RN(n6637), .QN(n5107) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][19]  ( .D(n6969), .E(
        n6814), .C(n1107), .RN(n6637), .QN(n5261) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][20]  ( .D(n6971), .E(
        n6814), .C(n1107), .RN(n6637), .QN(n5219) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][21]  ( .D(n6973), .E(
        n6814), .C(n1107), .RN(n6637), .QN(n5163) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][22]  ( .D(
        write_data_reg[22]), .E(n6814), .C(n1107), .RN(n6637), .QN(n5095) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][23]  ( .D(n6977), .E(
        n6814), .C(n1107), .RN(n6637), .QN(n5231) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][24]  ( .D(
        write_data_reg[24]), .E(n6814), .C(n1107), .RN(n6637), .QN(n5185) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][25]  ( .D(n6981), .E(
        n6813), .C(n1107), .RN(n6637), .QN(n5131) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][26]  ( .D(n6983), .E(
        n6813), .C(n1107), .RN(n6637), .QN(n5059) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][27]  ( .D(n6985), .E(
        n6813), .C(n1107), .RN(n6638), .QN(n5175) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][28]  ( .D(n6987), .E(
        n6813), .C(n1107), .RN(n6638), .QN(n5119) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][29]  ( .D(n6989), .E(
        n6813), .C(n1107), .RN(n6638), .QN(n5043) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][30]  ( .D(n6991), .E(
        n6813), .C(n1107), .RN(n6638), .QN(n4993) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[26][31]  ( .D(n6993), .E(
        n6813), .C(n1107), .RN(n6638), .QN(n5243) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][0]  ( .D(
        write_data_reg[0]), .E(n6892), .C(n1107), .RN(n6642), .QN(n4837) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][1]  ( .D(n6932), .E(
        n6892), .C(n1107), .RN(n6642), .QN(n5309) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][2]  ( .D(n6934), .E(
        n6892), .C(n1107), .RN(n6642), .QN(n4869) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][3]  ( .D(n6937), .E(
        n6892), .C(n1107), .RN(n6642), .QN(n4925) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][4]  ( .D(
        write_data_reg[4]), .E(n6891), .C(n1107), .RN(n6642), .QN(n4909) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][5]  ( .D(
        write_data_reg[5]), .E(n6891), .C(n1107), .RN(n6642), .QN(n4887) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][6]  ( .D(n6943), .E(
        n6891), .C(n1107), .RN(n6642), .QN(n4867) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][7]  ( .D(
        write_data_reg[7]), .E(n6891), .C(n1107), .RN(n6642), .QN(n4917) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][8]  ( .D(
        write_data_reg[8]), .E(n6891), .C(n1107), .RN(n6643), .QN(n4897) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][9]  ( .D(n6949), .E(
        n6891), .C(n1107), .RN(n6643), .QN(n4873) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][10]  ( .D(n6951), .E(
        n6891), .C(n1107), .RN(n6643), .QN(n4855) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][11]  ( .D(n6953), .E(
        n6890), .C(n1107), .RN(n6643), .QN(n4893) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][12]  ( .D(n6955), .E(
        n6890), .C(n1107), .RN(n6643), .QN(n4875) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][13]  ( .D(
        write_data_reg[13]), .E(n6890), .C(n1107), .RN(n6643), .QN(n4857) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][14]  ( .D(n6959), .E(
        n6890), .C(n1107), .RN(n6643), .QN(n5347) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][15]  ( .D(
        write_data_reg[15]), .E(n6890), .C(n1107), .RN(n6643), .QN(n4903) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][16]  ( .D(
        write_data_reg[16]), .E(n6890), .C(n1107), .RN(n6643), .QN(n4881) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][17]  ( .D(n6965), .E(
        n6890), .C(n1107), .RN(n6644), .QN(n4861) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][18]  ( .D(n6967), .E(
        n6889), .C(n1107), .RN(n6644), .QN(n4847) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][19]  ( .D(n6969), .E(
        n6889), .C(n1107), .RN(n6644), .QN(n4901) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][20]  ( .D(n6971), .E(
        n6889), .C(n1107), .RN(n6644), .QN(n4879) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][21]  ( .D(n6973), .E(
        n6889), .C(n1107), .RN(n6644), .QN(n4859) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][22]  ( .D(n6975), .E(
        n6889), .C(n1107), .RN(n6644), .QN(n4845) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][24]  ( .D(
        write_data_reg[24]), .E(n6889), .C(n1107), .RN(n6644), .QN(n4865) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][25]  ( .D(n6981), .E(
        n6889), .C(n1107), .RN(n6644), .QN(n4851) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][26]  ( .D(n6983), .E(
        n6888), .C(n1107), .RN(n6644), .QN(n4843) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][27]  ( .D(n6985), .E(
        n6888), .C(n1107), .RN(n6645), .QN(n4863) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][28]  ( .D(n6987), .E(
        n6888), .C(n1107), .RN(n6645), .QN(n4849) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][29]  ( .D(n6989), .E(
        n6888), .C(n1107), .RN(n6645), .QN(n4841) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][30]  ( .D(n6991), .E(
        n6888), .C(n1107), .RN(n6645), .QN(n4839) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[14][31]  ( .D(n6993), .E(
        n6888), .C(n1107), .RN(n6645), .QN(n4889) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][0]  ( .D(n6930), .E(
        n6912), .C(n1107), .RN(n6645), .QN(n4951) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][1]  ( .D(n6932), .E(
        n6912), .C(n1107), .RN(n6645), .QN(n5295) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][2]  ( .D(n6934), .E(
        n6912), .C(n1107), .RN(n6645), .QN(n5037) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][3]  ( .D(n6937), .E(
        n6912), .C(n1107), .RN(n6645), .QN(n5215) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][4]  ( .D(n6939), .E(
        n6911), .C(n1107), .RN(n6646), .QN(n5159) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][5]  ( .D(
        write_data_reg[5]), .E(n6911), .C(n1107), .RN(n6646), .QN(n5089) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][6]  ( .D(n6943), .E(
        n6911), .C(n1107), .RN(n6646), .QN(n5031) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][7]  ( .D(
        write_data_reg[7]), .E(n6911), .C(n1107), .RN(n6646), .QN(n5179) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][8]  ( .D(
        write_data_reg[8]), .E(n6911), .C(n1107), .RN(n6646), .QN(n5125) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][9]  ( .D(n6949), .E(
        n6911), .C(n1107), .RN(n6646), .QN(n5049) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][10]  ( .D(n6951), .E(
        n6911), .C(n1107), .RN(n6646), .QN(n4999) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][11]  ( .D(n6953), .E(
        n6910), .C(n1107), .RN(n6646), .QN(n5113) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][12]  ( .D(n6955), .E(
        n6910), .C(n1107), .RN(n6646), .QN(n5053) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][13]  ( .D(n6957), .E(
        n6910), .C(n1107), .RN(n6647), .QN(n5003) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][14]  ( .D(n6959), .E(
        n6910), .C(n1107), .RN(n6647), .QN(n4971) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][15]  ( .D(n6961), .E(
        n6910), .C(n1107), .RN(n6647), .QN(n5141) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][16]  ( .D(
        write_data_reg[16]), .E(n6910), .C(n1107), .RN(n6647), .QN(n5071) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][17]  ( .D(n6965), .E(
        n6910), .C(n1107), .RN(n6647), .QN(n5013) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][18]  ( .D(n6967), .E(
        n6909), .C(n1107), .RN(n6647), .QN(n4979) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][19]  ( .D(n6969), .E(
        n6909), .C(n1107), .RN(n6647), .QN(n5135) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][20]  ( .D(n6971), .E(
        n6909), .C(n1107), .RN(n6647), .QN(n5065) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][21]  ( .D(n6973), .E(
        n6909), .C(n1107), .RN(n6647), .QN(n5009) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][22]  ( .D(n6975), .E(
        n6909), .C(n1107), .RN(n6648), .QN(n4975) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][23]  ( .D(n6977), .E(
        n6909), .C(n1107), .RN(n6648), .QN(n5077) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][24]  ( .D(
        write_data_reg[24]), .E(n6909), .C(n1107), .RN(n6648), .QN(n5025) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][25]  ( .D(n6981), .E(
        n6908), .C(n1107), .RN(n6648), .QN(n4989) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][26]  ( .D(n6983), .E(
        n6908), .C(n1107), .RN(n6648), .QN(n4967) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][27]  ( .D(n6985), .E(
        n6908), .C(n1107), .RN(n6648), .QN(n5019) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][28]  ( .D(n6987), .E(
        n6908), .C(n1107), .RN(n6648), .QN(n4985) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][29]  ( .D(n6989), .E(
        n6908), .C(n1107), .RN(n6648), .QN(n4961) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][30]  ( .D(n6991), .E(
        n6908), .C(n1107), .RN(n6648), .QN(n4955) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[10][31]  ( .D(n6993), .E(
        n6908), .C(n1107), .RN(n6649), .QN(n5101) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][0]  ( .D(n6930), .E(n6777), .C(n1107), .RN(n6649), .QN(n4709) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][1]  ( .D(n6932), .E(n6777), .C(n1107), .RN(n6649), .QN(n4665) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][2]  ( .D(n6934), .E(n6777), .C(n1107), .RN(n6649), .QN(n4661) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][3]  ( .D(n6937), .E(n6777), .C(n1107), .RN(n6649), .QN(n4657) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][4]  ( .D(n6939), .E(n6776), .C(n1107), .RN(n6649), .QN(n4653) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][5]  ( .D(
        write_data_reg[5]), .E(n6776), .C(n1107), .RN(n6649), .QN(n4649) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][6]  ( .D(n6943), .E(n6776), .C(n1107), .RN(n6649), .QN(n4645) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][7]  ( .D(
        write_data_reg[7]), .E(n6776), .C(n1107), .RN(n6649), .QN(n4641) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][8]  ( .D(
        write_data_reg[8]), .E(n6776), .C(n1107), .RN(n6650), .QN(n4637) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][9]  ( .D(n6949), .E(n6776), .C(n1107), .RN(n6650), .QN(n4633) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][10]  ( .D(n6951), .E(
        n6776), .C(n1107), .RN(n6650), .QN(n4705) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][12]  ( .D(n6955), .E(
        n6775), .C(n1107), .RN(n6650), .QN(n4697) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][13]  ( .D(n6957), .E(
        n6775), .C(n1107), .RN(n6650), .QN(n4693) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][14]  ( .D(n6959), .E(
        n6775), .C(n1107), .RN(n6650), .QN(n4689) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][15]  ( .D(n6961), .E(
        n6775), .C(n1107), .RN(n6650), .QN(n4685) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][16]  ( .D(
        write_data_reg[16]), .E(n6775), .C(n1107), .RN(n6650), .QN(n4681) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][17]  ( .D(n6965), .E(
        n6775), .C(n1107), .RN(n6651), .QN(n4677) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][18]  ( .D(n6967), .E(
        n6774), .C(n1107), .RN(n6651), .QN(n4673) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][19]  ( .D(n6969), .E(
        n6774), .C(n1107), .RN(n6651), .QN(n4669) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][20]  ( .D(n6971), .E(
        n6774), .C(n1107), .RN(n6651), .QN(n4629) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][21]  ( .D(n6973), .E(
        n6774), .C(n1107), .RN(n6651), .QN(n4625) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][22]  ( .D(n6975), .E(
        n6774), .C(n1107), .RN(n6651), .QN(n4621) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][23]  ( .D(n6977), .E(
        n6774), .C(n1107), .RN(n6651), .QN(n4617) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][24]  ( .D(
        write_data_reg[24]), .E(n6774), .C(n1107), .RN(n6651), .QN(n4613) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][25]  ( .D(n6981), .E(
        n6773), .C(n1107), .RN(n6651), .QN(n4609) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][26]  ( .D(n6983), .E(
        n6773), .C(n1107), .RN(n6652), .QN(n4605) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][28]  ( .D(n6987), .E(
        n6773), .C(n1107), .RN(n6652), .QN(n4597) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][29]  ( .D(n6989), .E(
        n6773), .C(n1107), .RN(n6652), .QN(n4593) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][30]  ( .D(n6991), .E(
        n6773), .C(n1107), .RN(n6652), .QN(n4589) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][31]  ( .D(n6993), .E(
        n6773), .C(n1107), .RN(n6652), .QN(n4585) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][0]  ( .D(n6930), .E(
        n6852), .C(n1107), .RN(n6670), .QN(n4830) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][1]  ( .D(
        write_data_reg[1]), .E(n6852), .C(n1107), .RN(n6670), .QN(n5306) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][2]  ( .D(n6934), .E(
        n6852), .C(n1107), .RN(n6670), .QN(n4770) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][3]  ( .D(n6936), .E(
        n6852), .C(n1107), .RN(n6670), .QN(n4826) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][4]  ( .D(n6939), .E(
        n6851), .C(n1107), .RN(n6670), .QN(n4818) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][5]  ( .D(n6941), .E(
        n6851), .C(n1107), .RN(n6670), .QN(n4794) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][6]  ( .D(n6943), .E(
        n6851), .C(n1107), .RN(n6670), .QN(n4766) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][8]  ( .D(n6947), .E(
        n6851), .C(n1107), .RN(n6670), .QN(n4806) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][9]  ( .D(n6949), .E(
        n6851), .C(n1107), .RN(n6671), .QN(n4774) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][10]  ( .D(
        write_data_reg[10]), .E(n6851), .C(n1107), .RN(n6671), .QN(n4742) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][13]  ( .D(n6957), .E(
        n6850), .C(n1107), .RN(n6671), .QN(n4746) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][14]  ( .D(n6959), .E(
        n6850), .C(n1107), .RN(n6671), .QN(n4722) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][16]  ( .D(n6963), .E(
        n6850), .C(n1107), .RN(n6671), .QN(n4786) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][17]  ( .D(
        write_data_reg[17]), .E(n6850), .C(n1107), .RN(n6671), .QN(n4754) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][18]  ( .D(n6967), .E(
        n6849), .C(n1107), .RN(n6672), .QN(n4730) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][19]  ( .D(
        write_data_reg[19]), .E(n6849), .C(n1107), .RN(n6672), .QN(n4810) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][20]  ( .D(
        write_data_reg[20]), .E(n6849), .C(n1107), .RN(n6672), .QN(n4782) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][21]  ( .D(
        write_data_reg[21]), .E(n6849), .C(n1107), .RN(n6672), .QN(n4750) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][22]  ( .D(n6975), .E(
        n6849), .C(n1107), .RN(n6672), .QN(n4726) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][23]  ( .D(n6977), .E(
        n6849), .C(n1107), .RN(n6672), .QN(n4790) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][24]  ( .D(n6979), .E(
        n6849), .C(n1107), .RN(n6672), .QN(n4762) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][25]  ( .D(n6981), .E(
        n6848), .C(n1107), .RN(n6672), .QN(n4738) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][26]  ( .D(
        write_data_reg[26]), .E(n6848), .C(n1107), .RN(n6672), .QN(n4718) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][27]  ( .D(n6985), .E(
        n6848), .C(n1107), .RN(n6673), .QN(n4758) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][28]  ( .D(n6987), .E(
        n6848), .C(n1107), .RN(n6673), .QN(n4734) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][29]  ( .D(n6989), .E(
        n6848), .C(n1107), .RN(n6673), .QN(n4714) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][30]  ( .D(n6991), .E(
        n6848), .C(n1107), .RN(n6673), .QN(n4710) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[17][31]  ( .D(
        write_data_reg[31]), .E(n6848), .C(n1107), .RN(n6673), .QN(n4798) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[2][27]  ( .D(n6985), .E(
        n6773), .C(n1107), .RN(n6719), .QN(n4601) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][0]  ( .D(
        write_data_reg[0]), .E(n6787), .C(n1107), .RN(n6709), .Q(n5356) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][1]  ( .D(
        write_data_reg[1]), .E(n6787), .C(n1107), .RN(n6709), .Q(n5440) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][2]  ( .D(
        write_data_reg[2]), .E(n6787), .C(n1107), .RN(n6710), .Q(n5524) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][3]  ( .D(n6936), .E(n6787), .C(n1107), .RN(n6710), .Q(n5548) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][4]  ( .D(n6939), .E(n6786), .C(n1107), .RN(n6710), .Q(n5556) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][5]  ( .D(n6941), .E(n6786), .C(n1107), .RN(n6710), .Q(n5564) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][6]  ( .D(n6943), .E(n6786), .C(n1107), .RN(n6710), .Q(n5572) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][7]  ( .D(n6945), .E(n6786), .C(n1107), .RN(n6710), .Q(n5580) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][8]  ( .D(n6947), .E(n6786), .C(n1107), .RN(n6710), .Q(n5588) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][9]  ( .D(n6949), .E(n6786), .C(n1107), .RN(n6710), .Q(n5596) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][10]  ( .D(
        write_data_reg[10]), .E(n6786), .C(n1107), .RN(n6710), .Q(n5360) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][12]  ( .D(
        write_data_reg[12]), .E(n6785), .C(n1107), .RN(n6711), .Q(n5376) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][13]  ( .D(n6957), .E(
        n6785), .C(n1107), .RN(n6711), .Q(n5384) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][14]  ( .D(
        write_data_reg[14]), .E(n6785), .C(n1107), .RN(n6711), .Q(n5392) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][15]  ( .D(n6961), .E(
        n6785), .C(n1107), .RN(n6711), .Q(n5400) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][16]  ( .D(n6963), .E(
        n6785), .C(n1107), .RN(n6711), .Q(n5408) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][17]  ( .D(
        write_data_reg[17]), .E(n6785), .C(n1107), .RN(n6711), .Q(n5416) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][19]  ( .D(
        write_data_reg[19]), .E(n6784), .C(n1107), .RN(n6711), .Q(n5432) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][20]  ( .D(
        write_data_reg[20]), .E(n6784), .C(n1107), .RN(n6712), .Q(n5444) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][21]  ( .D(
        write_data_reg[21]), .E(n6784), .C(n1107), .RN(n6712), .Q(n5452) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][22]  ( .D(n6975), .E(
        n6784), .C(n1107), .RN(n6712), .Q(n5460) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][23]  ( .D(
        write_data_reg[23]), .E(n6784), .C(n1107), .RN(n6712), .Q(n5468) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][24]  ( .D(n6979), .E(
        n6784), .C(n1107), .RN(n6712), .Q(n5476) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][25]  ( .D(n6981), .E(
        n6783), .C(n1107), .RN(n6712), .Q(n5484) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][26]  ( .D(
        write_data_reg[26]), .E(n6783), .C(n1107), .RN(n6712), .Q(n5492) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][28]  ( .D(n6987), .E(
        n6783), .C(n1107), .RN(n6712), .Q(n5508) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][29]  ( .D(n6989), .E(
        n6783), .C(n1107), .RN(n6712), .Q(n5516) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][30]  ( .D(n6991), .E(
        n6783), .C(n1107), .RN(n6713), .Q(n5532) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][31]  ( .D(
        write_data_reg[31]), .E(n6783), .C(n1107), .RN(n6713), .Q(n5540) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][27]  ( .D(n6985), .E(
        n6783), .C(n1107), .RN(n6723), .Q(n5500) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][0]  ( .D(
        write_data_reg[0]), .E(n6802), .C(n1107), .RN(n6704), .Q(n5359) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][1]  ( .D(n6932), .E(n6802), .C(n1107), .RN(n6704), .Q(n5443) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][2]  ( .D(n6934), .E(n6802), .C(n1107), .RN(n6704), .Q(n5527) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][4]  ( .D(n6939), .E(n6802), .C(n1107), .RN(n6704), .Q(n5559) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][5]  ( .D(n6941), .E(n6801), .C(n1107), .RN(n6705), .Q(n5567) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][6]  ( .D(n6943), .E(n6801), .C(n1107), .RN(n6705), .Q(n5575) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][8]  ( .D(n6947), .E(n6801), .C(n1107), .RN(n6705), .Q(n5591) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][9]  ( .D(n6949), .E(n6801), .C(n1107), .RN(n6705), .Q(n5599) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][10]  ( .D(
        write_data_reg[10]), .E(n6801), .C(n1107), .RN(n6705), .Q(n5363) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][13]  ( .D(n6957), .E(
        n6801), .C(n1107), .RN(n6705), .Q(n5387) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][14]  ( .D(
        write_data_reg[14]), .E(n6801), .C(n1107), .RN(n6705), .Q(n5395) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][16]  ( .D(n6963), .E(
        n6800), .C(n1107), .RN(n6705), .Q(n5411) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][17]  ( .D(
        write_data_reg[17]), .E(n6800), .C(n1107), .RN(n6705), .Q(n5419) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][21]  ( .D(
        write_data_reg[21]), .E(n6800), .C(n1107), .RN(n6706), .Q(n5455) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][22]  ( .D(n6975), .E(
        n6800), .C(n1107), .RN(n6706), .Q(n5463) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][25]  ( .D(n6981), .E(
        n6800), .C(n1107), .RN(n6706), .Q(n5487) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][26]  ( .D(
        write_data_reg[26]), .E(n6800), .C(n1107), .RN(n6706), .Q(n5495) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][30]  ( .D(n6991), .E(
        n6799), .C(n1107), .RN(n6706), .Q(n5535) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][31]  ( .D(
        write_data_reg[31]), .E(n6799), .C(n1107), .RN(n6706), .Q(n5543) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][3]  ( .D(n6936), .E(n6799), .C(n1107), .RN(n6721), .Q(n5551) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][7]  ( .D(n6945), .E(n6799), .C(n1107), .RN(n6721), .Q(n5583) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][11]  ( .D(n6953), .E(
        n6799), .C(n1107), .RN(n6721), .Q(n5371) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][12]  ( .D(
        write_data_reg[12]), .E(n6799), .C(n1107), .RN(n6721), .Q(n5379) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][15]  ( .D(n6961), .E(
        n6799), .C(n1107), .RN(n6721), .Q(n5403) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][19]  ( .D(
        write_data_reg[19]), .E(n6798), .C(n1107), .RN(n6721), .Q(n5435) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][20]  ( .D(
        write_data_reg[20]), .E(n6798), .C(n1107), .RN(n6721), .Q(n5447) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][23]  ( .D(
        write_data_reg[23]), .E(n6798), .C(n1107), .RN(n6721), .Q(n5471) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][24]  ( .D(n6979), .E(
        n6798), .C(n1107), .RN(n6722), .Q(n5479) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][27]  ( .D(n6985), .E(
        n6798), .C(n1107), .RN(n6722), .Q(n5503) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][28]  ( .D(n6987), .E(
        n6798), .C(n1107), .RN(n6722), .Q(n5511) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][29]  ( .D(n6989), .E(
        n6798), .C(n1107), .RN(n6722), .Q(n5519) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[4][18]  ( .D(n6967), .E(
        n6784), .C(n1107), .RN(n6711), .Q(n5424) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[7][18]  ( .D(n6967), .E(
        n6800), .C(n1107), .RN(n6706), .Q(n5427) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][23]  ( .D(
        write_data_reg[23]), .E(n6838), .C(n1107), .RN(n6725), .QN(n4930) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][14]  ( .D(
        write_data_reg[14]), .E(n6838), .C(n1107), .RN(n6725), .QN(n4884) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][0]  ( .D(n6930), .E(
        n6842), .C(n1107), .RN(n6652), .QN(n5330) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][1]  ( .D(n6932), .E(
        n6842), .C(n1107), .RN(n6652), .QN(n5304) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][2]  ( .D(n6934), .E(
        n6842), .C(n1107), .RN(n6652), .QN(n4920) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][3]  ( .D(n6937), .E(
        n6842), .C(n1107), .RN(n6652), .QN(n5320) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][4]  ( .D(n6939), .E(
        n6841), .C(n1107), .RN(n6653), .QN(n4944) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][5]  ( .D(
        write_data_reg[5]), .E(n6841), .C(n1107), .RN(n6653), .QN(n4932) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][6]  ( .D(n6943), .E(
        n6841), .C(n1107), .RN(n6653), .QN(n4918) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][7]  ( .D(n6945), .E(
        n6841), .C(n1107), .RN(n6653), .QN(n4946) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][8]  ( .D(
        write_data_reg[8]), .E(n6841), .C(n1107), .RN(n6653), .QN(n4938) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][9]  ( .D(n6949), .E(
        n6841), .C(n1107), .RN(n6653), .QN(n5318) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][10]  ( .D(n6951), .E(
        n6841), .C(n1107), .RN(n6653), .QN(n4904) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][11]  ( .D(n6953), .E(
        n6840), .C(n1107), .RN(n6653), .QN(n4936) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][12]  ( .D(n6955), .E(
        n6840), .C(n1107), .RN(n6653), .QN(n4922) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][15]  ( .D(n6961), .E(
        n6840), .C(n1107), .RN(n6654), .QN(n4942) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][16]  ( .D(
        write_data_reg[16]), .E(n6840), .C(n1107), .RN(n6654), .QN(n4928) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][17]  ( .D(n6965), .E(
        n6840), .C(n1107), .RN(n6654), .QN(n4912) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][18]  ( .D(n6967), .E(
        n6840), .C(n1107), .RN(n6654), .QN(n4890) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][19]  ( .D(n6969), .E(
        n6840), .C(n1107), .RN(n6654), .QN(n4940) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][20]  ( .D(n6971), .E(
        n6839), .C(n1107), .RN(n6654), .QN(n4926) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][21]  ( .D(n6973), .E(
        n6839), .C(n1107), .RN(n6654), .QN(n4910) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][22]  ( .D(n6975), .E(
        n6839), .C(n1107), .RN(n6654), .QN(n5328) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][24]  ( .D(
        write_data_reg[24]), .E(n6839), .C(n1107), .RN(n6654), .QN(n5324) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][25]  ( .D(n6981), .E(
        n6839), .C(n1107), .RN(n6655), .QN(n4898) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][26]  ( .D(n6983), .E(
        n6839), .C(n1107), .RN(n6655), .QN(n4876) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][27]  ( .D(n6985), .E(
        n6839), .C(n1107), .RN(n6655), .QN(n4914) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][28]  ( .D(n6987), .E(
        n6838), .C(n1107), .RN(n6655), .QN(n4894) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][29]  ( .D(n6989), .E(
        n6838), .C(n1107), .RN(n6655), .QN(n4870) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][30]  ( .D(n6991), .E(
        n6838), .C(n1107), .RN(n6655), .QN(n4852) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][31]  ( .D(n6993), .E(
        n6838), .C(n1107), .RN(n6655), .QN(n4934) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][0]  ( .D(n6930), .E(
        n6832), .C(n1107), .RN(n6655), .QN(n5286) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][1]  ( .D(n6932), .E(
        n6832), .C(n1107), .RN(n6655), .QN(n5298) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][3]  ( .D(n6937), .E(
        n6832), .C(n1107), .RN(n6656), .QN(n5280) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][4]  ( .D(n6939), .E(
        n6831), .C(n1107), .RN(n6656), .QN(n5270) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][5]  ( .D(
        write_data_reg[5]), .E(n6831), .C(n1107), .RN(n6656), .QN(n5234) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][6]  ( .D(n6943), .E(
        n6831), .C(n1107), .RN(n6656), .QN(n5188) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][7]  ( .D(n6945), .E(
        n6831), .C(n1107), .RN(n6656), .QN(n5274) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][8]  ( .D(
        write_data_reg[8]), .E(n6831), .C(n1107), .RN(n6656), .QN(n5252) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][9]  ( .D(n6949), .E(
        n6831), .C(n1107), .RN(n6656), .QN(n5200) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][10]  ( .D(n6951), .E(
        n6831), .C(n1107), .RN(n6656), .QN(n5144) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][11]  ( .D(n6953), .E(
        n6830), .C(n1107), .RN(n6657), .QN(n5246) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][12]  ( .D(n6955), .E(
        n6830), .C(n1107), .RN(n6657), .QN(n5206) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][13]  ( .D(n6957), .E(
        n6830), .C(n1107), .RN(n6657), .QN(n5150) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][14]  ( .D(n6959), .E(
        n6830), .C(n1107), .RN(n6657), .QN(n5080) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][15]  ( .D(n6961), .E(
        n6830), .C(n1107), .RN(n6657), .QN(n5264) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][16]  ( .D(n6963), .E(
        n6830), .C(n1107), .RN(n6657), .QN(n5222) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][17]  ( .D(n6965), .E(
        n6830), .C(n1107), .RN(n6657), .QN(n5166) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][18]  ( .D(n6967), .E(
        n6829), .C(n1107), .RN(n6657), .QN(n5104) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][19]  ( .D(n6969), .E(
        n6829), .C(n1107), .RN(n6657), .QN(n5258) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][20]  ( .D(n6971), .E(
        n6829), .C(n1107), .RN(n6658), .QN(n5216) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][21]  ( .D(n6973), .E(
        n6829), .C(n1107), .RN(n6658), .QN(n5160) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][22]  ( .D(n6975), .E(
        n6829), .C(n1107), .RN(n6658), .QN(n5092) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][23]  ( .D(n6977), .E(
        n6829), .C(n1107), .RN(n6658), .QN(n5228) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][24]  ( .D(
        write_data_reg[24]), .E(n6829), .C(n1107), .RN(n6658), .QN(n5182) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][25]  ( .D(n6981), .E(
        n6828), .C(n1107), .RN(n6658), .QN(n5128) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][26]  ( .D(n6983), .E(
        n6828), .C(n1107), .RN(n6658), .QN(n5056) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][28]  ( .D(n6987), .E(
        n6828), .C(n1107), .RN(n6658), .QN(n5116) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][31]  ( .D(n6993), .E(
        n6828), .C(n1107), .RN(n6659), .QN(n5240) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][0]  ( .D(n6930), .E(
        n6822), .C(n1107), .RN(n6659), .QN(n5288) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][1]  ( .D(n6932), .E(
        n6822), .C(n1107), .RN(n6659), .QN(n5300) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][3]  ( .D(n6937), .E(
        n6822), .C(n1107), .RN(n6659), .QN(n5282) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][4]  ( .D(n6939), .E(
        n6821), .C(n1107), .RN(n6659), .QN(n5272) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][5]  ( .D(n6941), .E(
        n6821), .C(n1107), .RN(n6659), .QN(n5236) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][6]  ( .D(n6943), .E(
        n6821), .C(n1107), .RN(n6660), .QN(n5190) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][7]  ( .D(n6945), .E(
        n6821), .C(n1107), .RN(n6660), .QN(n5276) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][8]  ( .D(
        write_data_reg[8]), .E(n6821), .C(n1107), .RN(n6660), .QN(n5254) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][9]  ( .D(n6949), .E(
        n6821), .C(n1107), .RN(n6660), .QN(n5202) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][10]  ( .D(n6951), .E(
        n6821), .C(n1107), .RN(n6660), .QN(n5146) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][11]  ( .D(n6953), .E(
        n6820), .C(n1107), .RN(n6660), .QN(n5248) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][12]  ( .D(n6955), .E(
        n6820), .C(n1107), .RN(n6660), .QN(n5208) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][13]  ( .D(n6957), .E(
        n6820), .C(n1107), .RN(n6660), .QN(n5152) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][14]  ( .D(n6959), .E(
        n6820), .C(n1107), .RN(n6660), .QN(n5082) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][15]  ( .D(n6961), .E(
        n6820), .C(n1107), .RN(n6661), .QN(n5266) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][16]  ( .D(n6963), .E(
        n6820), .C(n1107), .RN(n6661), .QN(n5224) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][17]  ( .D(n6965), .E(
        n6820), .C(n1107), .RN(n6661), .QN(n5168) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][18]  ( .D(n6967), .E(
        n6819), .C(n1107), .RN(n6661), .QN(n5106) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][19]  ( .D(n6969), .E(
        n6819), .C(n1107), .RN(n6661), .QN(n5260) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][20]  ( .D(n6971), .E(
        n6819), .C(n1107), .RN(n6661), .QN(n5218) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][21]  ( .D(n6973), .E(
        n6819), .C(n1107), .RN(n6661), .QN(n5162) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][22]  ( .D(n6975), .E(
        n6819), .C(n1107), .RN(n6661), .QN(n5094) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][23]  ( .D(n6977), .E(
        n6819), .C(n1107), .RN(n6661), .QN(n5230) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][24]  ( .D(
        write_data_reg[24]), .E(n6819), .C(n1107), .RN(n6662), .QN(n5184) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][25]  ( .D(n6981), .E(
        n6818), .C(n1107), .RN(n6662), .QN(n5130) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][26]  ( .D(n6983), .E(
        n6818), .C(n1107), .RN(n6662), .QN(n5058) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][31]  ( .D(n6993), .E(
        n6818), .C(n1107), .RN(n6662), .QN(n5242) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][0]  ( .D(n6930), .E(
        n6812), .C(n1107), .RN(n6662), .QN(n5290) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][3]  ( .D(n6936), .E(
        n6812), .C(n1107), .RN(n6663), .QN(n5284) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][4]  ( .D(n6939), .E(
        n6811), .C(n1107), .RN(n6663), .QN(n5344) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][6]  ( .D(n6943), .E(
        n6811), .C(n1107), .RN(n6663), .QN(n5192) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][7]  ( .D(n6945), .E(
        n6811), .C(n1107), .RN(n6663), .QN(n5278) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][8]  ( .D(n6947), .E(
        n6811), .C(n1107), .RN(n6663), .QN(n5256) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][9]  ( .D(n6949), .E(
        n6811), .C(n1107), .RN(n6663), .QN(n5204) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][10]  ( .D(n6951), .E(
        n6811), .C(n1107), .RN(n6664), .QN(n5148) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][11]  ( .D(n6953), .E(
        n6810), .C(n1107), .RN(n6664), .QN(n5250) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][13]  ( .D(n6957), .E(
        n6810), .C(n1107), .RN(n6664), .QN(n5154) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][14]  ( .D(n6959), .E(
        n6810), .C(n1107), .RN(n6664), .QN(n5084) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][15]  ( .D(n6961), .E(
        n6810), .C(n1107), .RN(n6664), .QN(n5268) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][16]  ( .D(n6963), .E(
        n6810), .C(n1107), .RN(n6664), .QN(n5226) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][17]  ( .D(
        write_data_reg[17]), .E(n6810), .C(n1107), .RN(n6664), .QN(n5170) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][18]  ( .D(n6967), .E(
        n6809), .C(n1107), .RN(n6664), .QN(n5108) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][19]  ( .D(
        write_data_reg[19]), .E(n6809), .C(n1107), .RN(n6665), .QN(n5262) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][20]  ( .D(
        write_data_reg[20]), .E(n6809), .C(n1107), .RN(n6665), .QN(n5220) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][22]  ( .D(n6975), .E(
        n6809), .C(n1107), .RN(n6665), .QN(n5096) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][23]  ( .D(n6977), .E(
        n6809), .C(n1107), .RN(n6665), .QN(n5232) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][24]  ( .D(n6979), .E(
        n6809), .C(n1107), .RN(n6665), .QN(n5186) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][25]  ( .D(n6981), .E(
        n6808), .C(n1107), .RN(n6665), .QN(n5342) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][0]  ( .D(n6930), .E(
        n6897), .C(n1107), .RN(n6673), .QN(n4836) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][1]  ( .D(
        write_data_reg[1]), .E(n6897), .C(n1107), .RN(n6673), .QN(n5308) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][3]  ( .D(n6936), .E(
        n6897), .C(n1107), .RN(n6673), .QN(n4924) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][4]  ( .D(
        write_data_reg[4]), .E(n6896), .C(n1107), .RN(n6674), .QN(n4908) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][5]  ( .D(n6941), .E(
        n6896), .C(n1107), .RN(n6674), .QN(n4886) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][6]  ( .D(n6943), .E(
        n6896), .C(n1107), .RN(n6674), .QN(n4866) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][7]  ( .D(n6945), .E(
        n6896), .C(n1107), .RN(n6674), .QN(n4916) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][8]  ( .D(n6947), .E(
        n6896), .C(n1107), .RN(n6674), .QN(n4896) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][9]  ( .D(n6949), .E(
        n6896), .C(n1107), .RN(n6674), .QN(n4872) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][10]  ( .D(
        write_data_reg[10]), .E(n6896), .C(n1107), .RN(n6674), .QN(n4854) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][11]  ( .D(n6953), .E(
        n6895), .C(n1107), .RN(n6674), .QN(n4892) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][12]  ( .D(
        write_data_reg[12]), .E(n6895), .C(n1107), .RN(n6674), .QN(n4874) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][13]  ( .D(n6957), .E(
        n6895), .C(n1107), .RN(n6675), .QN(n4856) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][14]  ( .D(n6959), .E(
        n6895), .C(n1107), .RN(n6675), .QN(n5346) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][15]  ( .D(n6961), .E(
        n6895), .C(n1107), .RN(n6675), .QN(n4902) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][16]  ( .D(n6963), .E(
        n6895), .C(n1107), .RN(n6675), .QN(n4880) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][17]  ( .D(
        write_data_reg[17]), .E(n6895), .C(n1107), .RN(n6675), .QN(n4860) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][18]  ( .D(n6967), .E(
        n6894), .C(n1107), .RN(n6675), .QN(n4846) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][19]  ( .D(
        write_data_reg[19]), .E(n6894), .C(n1107), .RN(n6675), .QN(n4900) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][20]  ( .D(
        write_data_reg[20]), .E(n6894), .C(n1107), .RN(n6675), .QN(n4878) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][21]  ( .D(
        write_data_reg[21]), .E(n6894), .C(n1107), .RN(n6675), .QN(n4858) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][22]  ( .D(n6975), .E(
        n6894), .C(n1107), .RN(n6676), .QN(n4844) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][23]  ( .D(n6977), .E(
        n6894), .C(n1107), .RN(n6676), .QN(n4882) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][24]  ( .D(n6979), .E(
        n6894), .C(n1107), .RN(n6676), .QN(n4864) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][25]  ( .D(n6981), .E(
        n6893), .C(n1107), .RN(n6676), .QN(n4850) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][26]  ( .D(
        write_data_reg[26]), .E(n6893), .C(n1107), .RN(n6676), .QN(n4842) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][27]  ( .D(n6985), .E(
        n6893), .C(n1107), .RN(n6676), .QN(n4862) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][28]  ( .D(n6987), .E(
        n6893), .C(n1107), .RN(n6676), .QN(n4848) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][30]  ( .D(n6991), .E(
        n6893), .C(n1107), .RN(n6676), .QN(n4838) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][31]  ( .D(
        write_data_reg[31]), .E(n6893), .C(n1107), .RN(n6677), .QN(n4888) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][3]  ( .D(n6936), .E(
        n6887), .C(n1107), .RN(n6677), .QN(n5212) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][4]  ( .D(n6939), .E(
        n6887), .C(n1107), .RN(n6677), .QN(n5156) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][5]  ( .D(n6941), .E(
        n6887), .C(n1107), .RN(n6677), .QN(n5086) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][6]  ( .D(n6943), .E(
        n6887), .C(n1107), .RN(n6677), .QN(n5028) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][7]  ( .D(n6945), .E(
        n6886), .C(n1107), .RN(n6677), .QN(n5176) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][8]  ( .D(n6947), .E(
        n6886), .C(n1107), .RN(n6677), .QN(n5122) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][9]  ( .D(n6949), .E(
        n6886), .C(n1107), .RN(n6677), .QN(n5046) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][10]  ( .D(
        write_data_reg[10]), .E(n6886), .C(n1107), .RN(n6677), .QN(n4996) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][11]  ( .D(n6953), .E(
        n6886), .C(n1107), .RN(n6678), .QN(n5110) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][12]  ( .D(
        write_data_reg[12]), .E(n6886), .C(n1107), .RN(n6678), .QN(n5050) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][13]  ( .D(n6957), .E(
        n6886), .C(n1107), .RN(n6678), .QN(n5000) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][14]  ( .D(
        write_data_reg[14]), .E(n6885), .C(n1107), .RN(n6678), .QN(n4968) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][15]  ( .D(n6961), .E(
        n6885), .C(n1107), .RN(n6678), .QN(n5138) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][16]  ( .D(n6963), .E(
        n6885), .C(n1107), .RN(n6678), .QN(n5068) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][17]  ( .D(
        write_data_reg[17]), .E(n6885), .C(n1107), .RN(n6678), .QN(n5010) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][18]  ( .D(n6967), .E(
        n6885), .C(n1107), .RN(n6678), .QN(n4976) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][19]  ( .D(
        write_data_reg[19]), .E(n6885), .C(n1107), .RN(n6678), .QN(n5132) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][20]  ( .D(
        write_data_reg[20]), .E(n6885), .C(n1107), .RN(n6679), .QN(n5062) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][21]  ( .D(
        write_data_reg[21]), .E(n6884), .C(n1107), .RN(n6679), .QN(n5006) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][22]  ( .D(n6975), .E(
        n6884), .C(n1107), .RN(n6679), .QN(n4972) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][23]  ( .D(
        write_data_reg[23]), .E(n6884), .C(n1107), .RN(n6679), .QN(n5074) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][24]  ( .D(n6979), .E(
        n6884), .C(n1107), .RN(n6679), .QN(n5022) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][25]  ( .D(n6981), .E(
        n6884), .C(n1107), .RN(n6679), .QN(n4986) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][26]  ( .D(
        write_data_reg[26]), .E(n6884), .C(n1107), .RN(n6679), .QN(n4964) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][27]  ( .D(n6985), .E(
        n6884), .C(n1107), .RN(n6679), .QN(n5016) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][28]  ( .D(n6987), .E(
        n6883), .C(n1107), .RN(n6679), .QN(n4982) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][29]  ( .D(n6989), .E(
        n6883), .C(n1107), .RN(n6680), .QN(n4958) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][30]  ( .D(n6991), .E(
        n6883), .C(n1107), .RN(n6680), .QN(n4952) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][31]  ( .D(
        write_data_reg[31]), .E(n6883), .C(n1107), .RN(n6680), .QN(n5098) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][0]  ( .D(n6930), .E(
        n6917), .C(n1107), .RN(n6680), .QN(n4950) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][1]  ( .D(n6932), .E(
        n6917), .C(n1107), .RN(n6680), .QN(n5294) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][2]  ( .D(n6934), .E(
        n6917), .C(n1107), .RN(n6680), .QN(n5036) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][3]  ( .D(n6936), .E(
        n6917), .C(n1107), .RN(n6680), .QN(n5214) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][4]  ( .D(
        write_data_reg[4]), .E(n6916), .C(n1107), .RN(n6680), .QN(n5158) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][5]  ( .D(n6941), .E(
        n6916), .C(n1107), .RN(n6680), .QN(n5088) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][6]  ( .D(n6943), .E(
        n6916), .C(n1107), .RN(n6681), .QN(n5030) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][7]  ( .D(n6945), .E(
        n6916), .C(n1107), .RN(n6681), .QN(n5178) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][8]  ( .D(n6947), .E(
        n6916), .C(n1107), .RN(n6681), .QN(n5124) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][9]  ( .D(n6949), .E(
        n6916), .C(n1107), .RN(n6681), .QN(n5048) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][10]  ( .D(
        write_data_reg[10]), .E(n6916), .C(n1107), .RN(n6681), .QN(n4998) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][11]  ( .D(n6953), .E(
        n6915), .C(n1107), .RN(n6681), .QN(n5112) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][12]  ( .D(
        write_data_reg[12]), .E(n6915), .C(n1107), .RN(n6681), .QN(n5052) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][13]  ( .D(n6957), .E(
        n6915), .C(n1107), .RN(n6681), .QN(n5002) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][14]  ( .D(
        write_data_reg[14]), .E(n6915), .C(n1107), .RN(n6681), .QN(n4970) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][15]  ( .D(n6961), .E(
        n6915), .C(n1107), .RN(n6682), .QN(n5140) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][16]  ( .D(n6963), .E(
        n6915), .C(n1107), .RN(n6682), .QN(n5070) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][17]  ( .D(
        write_data_reg[17]), .E(n6915), .C(n1107), .RN(n6682), .QN(n5012) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][18]  ( .D(n6967), .E(
        n6914), .C(n1107), .RN(n6682), .QN(n4978) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][19]  ( .D(
        write_data_reg[19]), .E(n6914), .C(n1107), .RN(n6682), .QN(n5134) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][20]  ( .D(
        write_data_reg[20]), .E(n6914), .C(n1107), .RN(n6682), .QN(n5064) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][21]  ( .D(
        write_data_reg[21]), .E(n6914), .C(n1107), .RN(n6682), .QN(n5008) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][22]  ( .D(n6975), .E(
        n6914), .C(n1107), .RN(n6682), .QN(n4974) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][23]  ( .D(
        write_data_reg[23]), .E(n6914), .C(n1107), .RN(n6682), .QN(n5076) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][24]  ( .D(n6979), .E(
        n6914), .C(n1107), .RN(n6683), .QN(n5024) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][25]  ( .D(n6981), .E(
        n6913), .C(n1107), .RN(n6683), .QN(n4988) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][26]  ( .D(
        write_data_reg[26]), .E(n6913), .C(n1107), .RN(n6683), .QN(n4966) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][27]  ( .D(n6985), .E(
        n6913), .C(n1107), .RN(n6683), .QN(n5018) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][28]  ( .D(n6987), .E(
        n6913), .C(n1107), .RN(n6683), .QN(n4984) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][29]  ( .D(n6989), .E(
        n6913), .C(n1107), .RN(n6683), .QN(n4960) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][31]  ( .D(
        write_data_reg[31]), .E(n6913), .C(n1107), .RN(n6683), .QN(n5100) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][0]  ( .D(n6930), .E(n6907), .C(n1107), .RN(n6683), .QN(n5314) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][1]  ( .D(n6932), .E(n6907), .C(n1107), .RN(n6684), .QN(n5296) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][2]  ( .D(n6934), .E(n6907), .C(n1107), .RN(n6684), .QN(n5038) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][3]  ( .D(n6936), .E(n6907), .C(n1107), .RN(n6684), .QN(n5316) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][4]  ( .D(n6939), .E(n6906), .C(n1107), .RN(n6684), .QN(n5326) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][5]  ( .D(n6941), .E(n6906), .C(n1107), .RN(n6684), .QN(n5090) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][6]  ( .D(n6943), .E(n6906), .C(n1107), .RN(n6684), .QN(n5032) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][7]  ( .D(n6945), .E(n6906), .C(n1107), .RN(n6684), .QN(n5180) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][8]  ( .D(n6947), .E(n6906), .C(n1107), .RN(n6684), .QN(n5126) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][9]  ( .D(n6949), .E(n6906), .C(n1107), .RN(n6684), .QN(n5340) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][10]  ( .D(
        write_data_reg[10]), .E(n6906), .C(n1107), .RN(n6685), .QN(n5348) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][11]  ( .D(n6953), .E(
        n6905), .C(n1107), .RN(n6685), .QN(n5114) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][12]  ( .D(
        write_data_reg[12]), .E(n6905), .C(n1107), .RN(n6685), .QN(n5054) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][13]  ( .D(n6957), .E(
        n6905), .C(n1107), .RN(n6685), .QN(n5004) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][14]  ( .D(
        write_data_reg[14]), .E(n6905), .C(n1107), .RN(n6685), .QN(n5312) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][15]  ( .D(n6961), .E(
        n6905), .C(n1107), .RN(n6685), .QN(n5142) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][16]  ( .D(n6963), .E(
        n6905), .C(n1107), .RN(n6685), .QN(n5072) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][17]  ( .D(
        write_data_reg[17]), .E(n6905), .C(n1107), .RN(n6685), .QN(n5014) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][18]  ( .D(n6967), .E(
        n6904), .C(n1107), .RN(n6685), .QN(n4980) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][19]  ( .D(
        write_data_reg[19]), .E(n6904), .C(n1107), .RN(n6686), .QN(n5136) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][20]  ( .D(
        write_data_reg[20]), .E(n6904), .C(n1107), .RN(n6686), .QN(n5066) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][21]  ( .D(
        write_data_reg[21]), .E(n6904), .C(n1107), .RN(n6686), .QN(n5322) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][22]  ( .D(n6975), .E(
        n6904), .C(n1107), .RN(n6686), .QN(n5336) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][23]  ( .D(
        write_data_reg[23]), .E(n6904), .C(n1107), .RN(n6686), .QN(n5078) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][24]  ( .D(n6979), .E(
        n6904), .C(n1107), .RN(n6686), .QN(n5026) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][25]  ( .D(n6981), .E(
        n6903), .C(n1107), .RN(n6686), .QN(n5332) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][26]  ( .D(
        write_data_reg[26]), .E(n6903), .C(n1107), .RN(n6686), .QN(n5338) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][27]  ( .D(n6985), .E(
        n6903), .C(n1107), .RN(n6686), .QN(n5020) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][28]  ( .D(n6987), .E(
        n6903), .C(n1107), .RN(n6687), .QN(n5350) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][29]  ( .D(n6989), .E(
        n6903), .C(n1107), .RN(n6687), .QN(n4962) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[9][31]  ( .D(
        write_data_reg[31]), .E(n6903), .C(n1107), .RN(n6687), .QN(n5102) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][0]  ( .D(n6930), .E(n6782), .C(n1107), .RN(n6687), .QN(n4708) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][1]  ( .D(n6932), .E(n6782), .C(n1107), .RN(n6687), .QN(n4664) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][2]  ( .D(n6934), .E(n6782), .C(n1107), .RN(n6687), .QN(n4660) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][3]  ( .D(n6936), .E(n6782), .C(n1107), .RN(n6687), .QN(n4656) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][4]  ( .D(
        write_data_reg[4]), .E(n6781), .C(n1107), .RN(n6687), .QN(n4652) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][5]  ( .D(n6941), .E(n6781), .C(n1107), .RN(n6688), .QN(n4648) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][6]  ( .D(n6943), .E(n6781), .C(n1107), .RN(n6688), .QN(n4644) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][7]  ( .D(n6945), .E(n6781), .C(n1107), .RN(n6688), .QN(n4640) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][8]  ( .D(n6947), .E(n6781), .C(n1107), .RN(n6688), .QN(n4636) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][9]  ( .D(n6949), .E(n6781), .C(n1107), .RN(n6688), .QN(n4632) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][10]  ( .D(
        write_data_reg[10]), .E(n6781), .C(n1107), .RN(n6688), .QN(n4704) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][12]  ( .D(
        write_data_reg[12]), .E(n6780), .C(n1107), .RN(n6688), .QN(n4696) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][13]  ( .D(n6957), .E(
        n6780), .C(n1107), .RN(n6688), .QN(n4692) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][14]  ( .D(
        write_data_reg[14]), .E(n6780), .C(n1107), .RN(n6688), .QN(n4688) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][15]  ( .D(n6961), .E(
        n6780), .C(n1107), .RN(n6689), .QN(n4684) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][16]  ( .D(n6963), .E(
        n6780), .C(n1107), .RN(n6689), .QN(n4680) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][17]  ( .D(
        write_data_reg[17]), .E(n6780), .C(n1107), .RN(n6689), .QN(n4676) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][18]  ( .D(n6967), .E(
        n6780), .C(n1107), .RN(n6689), .QN(n4672) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][19]  ( .D(
        write_data_reg[19]), .E(n6779), .C(n1107), .RN(n6689), .QN(n4668) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][20]  ( .D(
        write_data_reg[20]), .E(n6779), .C(n1107), .RN(n6689), .QN(n4628) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][21]  ( .D(
        write_data_reg[21]), .E(n6779), .C(n1107), .RN(n6689), .QN(n4624) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][22]  ( .D(n6975), .E(
        n6779), .C(n1107), .RN(n6689), .QN(n4620) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][24]  ( .D(n6979), .E(
        n6779), .C(n1107), .RN(n6689), .QN(n4612) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][25]  ( .D(n6981), .E(
        n6779), .C(n1107), .RN(n6690), .QN(n4608) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][26]  ( .D(
        write_data_reg[26]), .E(n6779), .C(n1107), .RN(n6690), .QN(n4604) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][29]  ( .D(n6989), .E(
        n6778), .C(n1107), .RN(n6690), .QN(n4592) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][30]  ( .D(n6991), .E(
        n6778), .C(n1107), .RN(n6690), .QN(n4588) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][31]  ( .D(
        write_data_reg[31]), .E(n6778), .C(n1107), .RN(n6690), .QN(n4584) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][0]  ( .D(n6930), .E(n6772), .C(n1107), .RN(n6690), .QN(n4706) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][1]  ( .D(n6932), .E(n6772), .C(n1107), .RN(n6690), .QN(n4662) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][2]  ( .D(n6934), .E(n6772), .C(n1107), .RN(n6690), .QN(n4658) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][3]  ( .D(n6936), .E(n6772), .C(n1107), .RN(n6690), .QN(n4654) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][4]  ( .D(n6939), .E(n6771), .C(n1107), .RN(n6691), .QN(n4650) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][5]  ( .D(n6941), .E(n6771), .C(n1107), .RN(n6691), .QN(n4646) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][6]  ( .D(n6943), .E(n6771), .C(n1107), .RN(n6691), .QN(n4642) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][7]  ( .D(n6945), .E(n6771), .C(n1107), .RN(n6691), .QN(n4638) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][8]  ( .D(n6947), .E(n6771), .C(n1107), .RN(n6691), .QN(n4634) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][9]  ( .D(n6949), .E(n6771), .C(n1107), .RN(n6691), .QN(n4630) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][10]  ( .D(
        write_data_reg[10]), .E(n6771), .C(n1107), .RN(n6691), .QN(n4702) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][11]  ( .D(n6953), .E(
        n6770), .C(n1107), .RN(n6691), .QN(n4698) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][12]  ( .D(
        write_data_reg[12]), .E(n6770), .C(n1107), .RN(n6691), .QN(n4694) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][13]  ( .D(n6957), .E(
        n6770), .C(n1107), .RN(n6692), .QN(n4690) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][14]  ( .D(
        write_data_reg[14]), .E(n6770), .C(n1107), .RN(n6692), .QN(n4686) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][15]  ( .D(n6961), .E(
        n6770), .C(n1107), .RN(n6692), .QN(n4682) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][16]  ( .D(n6963), .E(
        n6770), .C(n1107), .RN(n6692), .QN(n4678) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][17]  ( .D(
        write_data_reg[17]), .E(n6770), .C(n1107), .RN(n6692), .QN(n4674) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][18]  ( .D(n6967), .E(
        n6769), .C(n1107), .RN(n6692), .QN(n4670) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][19]  ( .D(
        write_data_reg[19]), .E(n6769), .C(n1107), .RN(n6692), .QN(n4666) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][20]  ( .D(
        write_data_reg[20]), .E(n6769), .C(n1107), .RN(n6692), .QN(n4626) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][21]  ( .D(
        write_data_reg[21]), .E(n6769), .C(n1107), .RN(n6692), .QN(n4622) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][22]  ( .D(n6975), .E(
        n6769), .C(n1107), .RN(n6693), .QN(n4618) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][23]  ( .D(
        write_data_reg[23]), .E(n6769), .C(n1107), .RN(n6693), .QN(n4614) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][24]  ( .D(n6979), .E(
        n6769), .C(n1107), .RN(n6693), .QN(n4610) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][25]  ( .D(n6981), .E(
        n6768), .C(n1107), .RN(n6693), .QN(n4606) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][26]  ( .D(
        write_data_reg[26]), .E(n6768), .C(n1107), .RN(n6693), .QN(n4602) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][28]  ( .D(n6987), .E(
        n6768), .C(n1107), .RN(n6693), .QN(n4594) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][29]  ( .D(n6989), .E(
        n6768), .C(n1107), .RN(n6693), .QN(n4590) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][30]  ( .D(n6991), .E(
        n6768), .C(n1107), .RN(n6693), .QN(n4586) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][31]  ( .D(
        write_data_reg[31]), .E(n6768), .C(n1107), .RN(n6693), .QN(n4582) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[31][13]  ( .D(n6957), .E(
        n6838), .C(n1107), .RN(n6694), .QN(n4906) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][0]  ( .D(n6930), .E(
        n6883), .C(n1107), .RN(n6694), .QN(n4948) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][1]  ( .D(n6932), .E(
        n6883), .C(n1107), .RN(n6694), .QN(n5292) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[13][2]  ( .D(n6934), .E(
        n6883), .C(n1107), .RN(n6694), .QN(n5034) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[22][0]  ( .D(
        write_data_reg[0]), .E(n6877), .C(n1107), .RN(n6713), .QN(n5692) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][11]  ( .D(n6953), .E(
        n6778), .C(n1107), .RN(n6720), .QN(n4700) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][23]  ( .D(
        write_data_reg[23]), .E(n6778), .C(n1107), .RN(n6720), .QN(n4616) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][27]  ( .D(n6985), .E(
        n6778), .C(n1107), .RN(n6720), .QN(n4600) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[3][28]  ( .D(n6987), .E(
        n6778), .C(n1107), .RN(n6720), .QN(n4596) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[1][27]  ( .D(n6985), .E(
        n6768), .C(n1107), .RN(n6720), .QN(n4598) );
  MUX22 \execute/alu/sll_175/M1_1_13  ( .A(\execute/alu/sll_175/ML_int[1][13] ), .B(\execute/alu/sll_175/ML_int[1][11] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][13] ) );
  MUX22 \execute/alu/sll_175/M1_1_7  ( .A(\execute/alu/sll_175/ML_int[1][7] ), 
        .B(\execute/alu/sll_175/ML_int[1][5] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][7] ) );
  MUX22 \execute/alu/sll_175/M1_4_24  ( .A(\execute/alu/sll_175/ML_int[4][24] ), .B(\execute/alu/sll_175/ML_int[4][8] ), .S(n6342), .Q(
        \execute/alu/sll_175/ML_int[5][24] ) );
  MUX22 \execute/alu/sll_175/M1_1_3  ( .A(\execute/alu/sll_175/ML_int[1][3] ), 
        .B(\execute/alu/sll_175/ML_int[1][1] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][3] ) );
  MUX22 \execute/alu/sll_175/M1_1_6  ( .A(\execute/alu/sll_175/ML_int[1][6] ), 
        .B(\execute/alu/sll_175/ML_int[1][4] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][6] ) );
  MUX22 \execute/alu/sll_175/M1_1_11  ( .A(\execute/alu/sll_175/ML_int[1][11] ), .B(\execute/alu/sll_175/ML_int[1][9] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][11] ) );
  MUX22 \execute/alu/sll_175/M1_1_5  ( .A(\execute/alu/sll_175/ML_int[1][5] ), 
        .B(\execute/alu/sll_175/ML_int[1][3] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][5] ) );
  MUX22 \execute/alu/sll_175/M1_1_4  ( .A(\execute/alu/sll_175/ML_int[1][4] ), 
        .B(\execute/alu/sll_175/ML_int[1][2] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][4] ) );
  MUX22 \execute/alu/sll_175/M1_3_23  ( .A(\execute/alu/sll_175/ML_int[3][23] ), .B(\execute/alu/sll_175/ML_int[3][15] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][23] ) );
  MUX22 \execute/alu/sll_175/M1_4_23  ( .A(\execute/alu/sll_175/ML_int[4][23] ), .B(n1211), .S(n6342), .Q(\execute/alu/sll_175/ML_int[5][23] ) );
  MUX22 \execute/alu/sll_175/M1_2_13  ( .A(\execute/alu/sll_175/ML_int[2][13] ), .B(\execute/alu/sll_175/ML_int[2][9] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][13] ) );
  MUX22 \execute/alu/sll_175/M1_2_17  ( .A(\execute/alu/sll_175/ML_int[2][17] ), .B(\execute/alu/sll_175/ML_int[2][13] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][17] ) );
  MUX22 \execute/alu/sll_175/M1_1_24  ( .A(\execute/alu/sll_175/ML_int[1][24] ), .B(\execute/alu/sll_175/ML_int[1][22] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][24] ) );
  MUX22 \execute/alu/sll_175/M1_1_22  ( .A(\execute/alu/sll_175/ML_int[1][22] ), .B(\execute/alu/sll_175/ML_int[1][20] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][22] ) );
  MUX22 \execute/alu/sll_175/M1_1_23  ( .A(\execute/alu/sll_175/ML_int[1][23] ), .B(\execute/alu/sll_175/ML_int[1][21] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][23] ) );
  MUX22 \execute/alu/sll_175/M1_0_19  ( .A(n1447), .B(n1445), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][19] ) );
  MUX22 \execute/alu/sll_175/M1_0_10  ( .A(n1428), .B(n1427), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][10] ) );
  MUX22 \execute/alu/sll_175/M1_2_7  ( .A(\execute/alu/sll_175/ML_int[2][7] ), 
        .B(\execute/alu/sll_175/ML_int[2][3] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][7] ) );
  MUX22 \execute/alu/sll_175/M1_2_14  ( .A(\execute/alu/sll_175/ML_int[2][14] ), .B(\execute/alu/sll_175/ML_int[2][10] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][14] ) );
  MUX22 \execute/alu/sll_175/M1_2_10  ( .A(\execute/alu/sll_175/ML_int[2][10] ), .B(\execute/alu/sll_175/ML_int[2][6] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][10] ) );
  MUX22 \execute/alu/sll_175/M1_1_2  ( .A(\execute/alu/sll_175/ML_int[1][2] ), 
        .B(n5812), .S(n5820), .Q(\execute/alu/sll_175/ML_int[2][2] ) );
  MUX22 \execute/alu/sll_175/M1_2_5  ( .A(\execute/alu/sll_175/ML_int[2][5] ), 
        .B(n5810), .S(n6758), .Q(\execute/alu/sll_175/ML_int[3][5] ) );
  MUX22 \execute/alu/sll_175/M1_2_15  ( .A(\execute/alu/sll_175/ML_int[2][15] ), .B(\execute/alu/sll_175/ML_int[2][11] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][15] ) );
  MUX22 \execute/alu/sll_175/M1_2_8  ( .A(\execute/alu/sll_175/ML_int[2][8] ), 
        .B(\execute/alu/sll_175/ML_int[2][4] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][8] ) );
  MUX22 \execute/alu/sll_175/M1_2_6  ( .A(\execute/alu/sll_175/ML_int[2][6] ), 
        .B(\execute/alu/sll_175/ML_int[2][2] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][6] ) );
  MUX22 \execute/alu/sll_175/M1_3_26  ( .A(\execute/alu/sll_175/ML_int[3][26] ), .B(\execute/alu/sll_175/ML_int[3][18] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][26] ) );
  MUX22 \execute/alu/sll_175/M1_4_26  ( .A(\execute/alu/sll_175/ML_int[4][26] ), .B(\execute/alu/sll_175/ML_int[4][10] ), .S(n6342), .Q(
        \execute/alu/sll_175/ML_int[5][26] ) );
  MUX22 \execute/alu/sll_175/M1_2_26  ( .A(\execute/alu/sll_175/ML_int[2][26] ), .B(\execute/alu/sll_175/ML_int[2][22] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][26] ) );
  MUX22 \execute/alu/sll_175/M1_1_9  ( .A(\execute/alu/sll_175/ML_int[1][9] ), 
        .B(\execute/alu/sll_175/ML_int[1][7] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][9] ) );
  MUX22 \execute/alu/sll_175/M1_3_30  ( .A(\execute/alu/sll_175/ML_int[3][30] ), .B(\execute/alu/sll_175/ML_int[3][22] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][30] ) );
  MUX22 \execute/alu/sll_175/M1_2_29  ( .A(\execute/alu/sll_175/ML_int[2][29] ), .B(\execute/alu/sll_175/ML_int[2][25] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][29] ) );
  MUX22 \execute/alu/sll_175/M1_3_29  ( .A(\execute/alu/sll_175/ML_int[3][29] ), .B(\execute/alu/sll_175/ML_int[3][21] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][29] ) );
  MUX22 \execute/alu/sll_175/M1_4_29  ( .A(\execute/alu/sll_175/ML_int[4][29] ), .B(\execute/alu/sll_175/ML_int[4][13] ), .S(n6342), .Q(
        \execute/alu/sll_175/ML_int[5][29] ) );
  MUX22 \execute/alu/sll_175/M1_2_25  ( .A(\execute/alu/sll_175/ML_int[2][25] ), .B(\execute/alu/sll_175/ML_int[2][21] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][25] ) );
  MUX22 \execute/alu/sll_175/M1_3_25  ( .A(\execute/alu/sll_175/ML_int[3][25] ), .B(\execute/alu/sll_175/ML_int[3][17] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][25] ) );
  MUX22 \execute/alu/sll_175/M1_4_25  ( .A(\execute/alu/sll_175/ML_int[4][25] ), .B(\execute/alu/sll_175/ML_int[4][9] ), .S(n6342), .Q(
        \execute/alu/sll_175/ML_int[5][25] ) );
  MUX22 \execute/alu/sll_175/M1_3_21  ( .A(\execute/alu/sll_175/ML_int[3][21] ), .B(\execute/alu/sll_175/ML_int[3][13] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][21] ) );
  MUX22 \execute/alu/sll_175/M1_4_17  ( .A(\execute/alu/sll_175/ML_int[4][17] ), .B(n5811), .S(n6343), .Q(\execute/alu/sll_175/ML_int[5][17] ) );
  MUX22 \execute/alu/sll_175/M1_3_28  ( .A(\execute/alu/sll_175/ML_int[3][28] ), .B(\execute/alu/sll_175/ML_int[3][20] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][28] ) );
  MUX22 \execute/alu/sll_175/M1_4_28  ( .A(\execute/alu/sll_175/ML_int[4][28] ), .B(\execute/alu/sll_175/ML_int[4][12] ), .S(n6342), .Q(
        \execute/alu/sll_175/ML_int[5][28] ) );
  MUX22 \execute/alu/sll_175/M1_3_27  ( .A(\execute/alu/sll_175/ML_int[3][27] ), .B(\execute/alu/sll_175/ML_int[3][19] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][27] ) );
  MUX22 \execute/alu/sll_175/M1_4_27  ( .A(\execute/alu/sll_175/ML_int[4][27] ), .B(\execute/alu/sll_175/ML_int[4][11] ), .S(n6342), .Q(
        \execute/alu/sll_175/ML_int[5][27] ) );
  MUX22 \execute/alu/sll_175/M1_2_24  ( .A(\execute/alu/sll_175/ML_int[2][24] ), .B(\execute/alu/sll_175/ML_int[2][20] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][24] ) );
  MUX22 \execute/alu/sll_175/M1_3_24  ( .A(\execute/alu/sll_175/ML_int[3][24] ), .B(\execute/alu/sll_175/ML_int[3][16] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][24] ) );
  MUX22 \execute/alu/sll_175/M1_3_8  ( .A(\execute/alu/sll_175/ML_int[3][8] ), 
        .B(n5808), .S(n5819), .Q(\execute/alu/sll_175/ML_int[4][8] ) );
  MUX22 \execute/alu/sll_175/M1_3_9  ( .A(\execute/alu/sll_175/ML_int[3][9] ), 
        .B(n1225), .S(n5819), .Q(\execute/alu/sll_175/ML_int[4][9] ) );
  MUX22 \execute/alu/sll_175/M1_3_14  ( .A(\execute/alu/sll_175/ML_int[3][14] ), .B(\execute/alu/sll_175/ML_int[3][6] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][14] ) );
  MUX22 \execute/alu/sll_175/M1_3_10  ( .A(\execute/alu/sll_175/ML_int[3][10] ), .B(n1218), .S(n5819), .Q(\execute/alu/sll_175/ML_int[4][10] ) );
  MUX22 \execute/alu/sll_175/M1_3_11  ( .A(\execute/alu/sll_175/ML_int[3][11] ), .B(n1224), .S(n5819), .Q(\execute/alu/sll_175/ML_int[4][11] ) );
  MUX22 \execute/alu/sll_175/M1_3_12  ( .A(\execute/alu/sll_175/ML_int[3][12] ), .B(\execute/alu/sll_175/ML_int[3][4] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][12] ) );
  MUX22 \execute/alu/sll_175/M1_2_23  ( .A(\execute/alu/sll_175/ML_int[2][23] ), .B(\execute/alu/sll_175/ML_int[2][19] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][23] ) );
  MUX22 \execute/alu/sll_175/M1_1_19  ( .A(\execute/alu/sll_175/ML_int[1][19] ), .B(\execute/alu/sll_175/ML_int[1][17] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][19] ) );
  DF1 \memory/read_data_reg[2]  ( .D(ram_word[2]), .C(clk), .QN(n5640) );
  DF1 \memory/read_data_reg[4]  ( .D(ram_word[4]), .C(clk), .QN(n5644) );
  DF1 \memory/read_data_reg[31]  ( .D(ram_word[31]), .C(clk), .QN(n5634) );
  DF1 \memory/read_data_reg[5]  ( .D(ram_word[5]), .C(clk), .QN(n5638) );
  DF1 \memory/read_data_reg[3]  ( .D(ram_word[3]), .C(clk), .QN(n5648) );
  DF1 \memory/address_WB_reg[2]  ( .D(ram_adr[2]), .C(clk), .QN(n5641) );
  DF1 \memory/address_WB_reg[31]  ( .D(ram_adr[31]), .C(clk), .QN(n5635) );
  DF1 \memory/address_WB_reg[5]  ( .D(ram_adr[5]), .C(clk), .QN(n5639) );
  DF1 \memory/address_WB_reg[3]  ( .D(ram_adr[3]), .C(clk), .QN(n5649) );
  DF1 \memory/read_data_reg[12]  ( .D(ram_word[12]), .C(clk), .QN(n5676) );
  DF1 \memory/read_data_reg[21]  ( .D(ram_word[21]), .C(clk), .QN(n5646) );
  DF1 \memory/read_data_reg[10]  ( .D(ram_word[10]), .C(clk), .QN(n5680) );
  DF1 \memory/read_data_reg[19]  ( .D(ram_word[19]), .C(clk), .QN(n5670) );
  DF1 \memory/read_data_reg[20]  ( .D(ram_word[20]), .C(clk), .QN(n5660) );
  DF1 \memory/read_data_reg[24]  ( .D(ram_word[24]), .C(clk), .QN(n5656) );
  DF1 \memory/read_data_reg[7]  ( .D(ram_word[7]), .C(clk), .QN(n5672) );
  DF1 \memory/read_data_reg[8]  ( .D(ram_word[8]), .C(clk), .QN(n5666) );
  DF1 \memory/read_data_reg[11]  ( .D(ram_word[11]), .C(clk), .QN(n5684) );
  DF1 \memory/read_data_reg[6]  ( .D(ram_word[6]), .C(clk), .QN(n5688) );
  DF1 \memory/read_data_reg[23]  ( .D(ram_word[23]), .C(clk), .QN(n5650) );
  DF1 \memory/read_data_reg[13]  ( .D(ram_word[13]), .C(clk), .QN(n5686) );
  DF1 \memory/read_data_reg[16]  ( .D(ram_word[16]), .C(clk), .QN(n5678) );
  DF1 \memory/read_data_reg[22]  ( .D(ram_word[22]), .C(clk), .QN(n5652) );
  DF1 \memory/read_data_reg[15]  ( .D(ram_word[15]), .C(clk), .QN(n5668) );
  DF1 \memory/read_data_reg[17]  ( .D(ram_word[17]), .C(clk), .QN(n5682) );
  DF1 \memory/read_data_reg[14]  ( .D(ram_word[14]), .C(clk), .QN(n5664) );
  DF1 \memory/read_data_reg[26]  ( .D(ram_word[26]), .C(clk), .QN(n5636) );
  DF1 \memory/read_data_reg[25]  ( .D(ram_word[25]), .C(clk), .QN(n5662) );
  DF1 \memory/read_data_reg[18]  ( .D(ram_word[18]), .C(clk), .QN(n5654) );
  DF1 \memory/read_data_reg[27]  ( .D(ram_word[27]), .C(clk), .QN(n5632) );
  DF1 \memory/address_WB_reg[12]  ( .D(ram_adr[12]), .C(clk), .QN(n5677) );
  DF1 \memory/address_WB_reg[19]  ( .D(ram_adr[19]), .C(clk), .QN(n5671) );
  DF1 \memory/address_WB_reg[24]  ( .D(ram_adr[24]), .C(clk), .QN(n5657) );
  DF1 \memory/address_WB_reg[7]  ( .D(ram_adr[7]), .C(clk), .QN(n5673) );
  DF1 \memory/address_WB_reg[8]  ( .D(ram_adr[8]), .C(clk), .QN(n5667) );
  DF1 \memory/address_WB_reg[11]  ( .D(ram_adr[11]), .C(clk), .QN(n5685) );
  DF1 \memory/address_WB_reg[6]  ( .D(ram_adr[6]), .C(clk), .QN(n5689) );
  DF1 \memory/address_WB_reg[23]  ( .D(ram_adr[23]), .C(clk), .QN(n5651) );
  DF1 \memory/address_WB_reg[13]  ( .D(ram_adr[13]), .C(clk), .QN(n5687) );
  DF1 \memory/address_WB_reg[22]  ( .D(ram_adr[22]), .C(clk), .QN(n5653) );
  DF1 \memory/address_WB_reg[15]  ( .D(ram_adr[15]), .C(clk), .QN(n5669) );
  DF1 \memory/address_WB_reg[14]  ( .D(ram_adr[14]), .C(clk), .QN(n5665) );
  DF1 \memory/address_WB_reg[26]  ( .D(ram_adr[26]), .C(clk), .QN(n5637) );
  DF1 \memory/address_WB_reg[25]  ( .D(ram_adr[25]), .C(clk), .QN(n5663) );
  DF1 \memory/address_WB_reg[18]  ( .D(ram_adr[18]), .C(clk), .QN(n5655) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[27][29]  ( .D(n6989), .E(
        n6818), .C(n1107), .RN(n6662), .QN(n5042) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[27][30]  ( .D(n6991), .E(
        n6818), .C(n1107), .RN(n6662), .QN(n4992) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[25][2]  ( .D(n6934), .E(
        n6812), .C(n1107), .RN(n6663), .QN(n5198) );
  DF1 \memory/read_data_reg[9]  ( .D(ram_word[9]), .C(clk), .QN(n5674) );
  DF1 \memory/read_data_reg[28]  ( .D(ram_word[28]), .C(clk), .QN(n5628) );
  DF1 \memory/read_data_reg[29]  ( .D(ram_word[29]), .C(clk), .QN(n5630) );
  DF1 \memory/read_data_reg[30]  ( .D(ram_word[30]), .C(clk), .QN(n5690) );
  DF1 \instruction_decode/imm_reg[0]  ( .D(inst_out[0]), .C(clk), .Q(n5946) );
  DF1 \memory/address_WB_reg[27]  ( .D(ram_adr[27]), .C(clk), .QN(n5633) );
  DF1 \memory/address_WB_reg[28]  ( .D(ram_adr[28]), .C(clk), .QN(n5629) );
  DF1 \memory/address_WB_reg[29]  ( .D(ram_adr[29]), .C(clk), .QN(n5631) );
  DF1 \memory/address_WB_reg[30]  ( .D(ram_adr[30]), .C(clk), .QN(n5691) );
  DF1 \memory/address_WB_reg[9]  ( .D(ram_adr[9]), .C(clk), .QN(n5675) );
  MUX21 \execute/alu/sll_175/M1_0_4  ( .A(n6347), .B(n6349), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][4] ) );
  MUX21 \execute/alu/sll_175/M1_0_12  ( .A(n6345), .B(n6344), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][12] ) );
  MUX21 \execute/alu/sll_175/M1_0_13  ( .A(n6346), .B(n6345), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][13] ) );
  MUX21 \execute/alu/sll_175/M1_0_5  ( .A(n1422), .B(n6347), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][5] ) );
  MUX21 \execute/alu/sll_175/M1_0_11  ( .A(n6344), .B(n1428), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][11] ) );
  MUX21 \execute/alu/sll_175/M1_0_16  ( .A(n6222), .B(n5829), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][16] ) );
  MUX21 \execute/alu/sll_175/M1_0_15  ( .A(n5829), .B(n5830), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][15] ) );
  MUX21 \execute/alu/sll_175/M1_0_14  ( .A(n5830), .B(n6346), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][14] ) );
  MUX21 \execute/alu/sll_175/M1_1_17  ( .A(\execute/alu/sll_175/ML_int[1][17] ), .B(\execute/alu/sll_175/ML_int[1][15] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][17] ) );
  MUX21 \execute/alu/sll_175/M1_1_18  ( .A(\execute/alu/sll_175/ML_int[1][18] ), .B(\execute/alu/sll_175/ML_int[1][16] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][18] ) );
  MUX21 \execute/alu/sll_175/M1_1_16  ( .A(\execute/alu/sll_175/ML_int[1][16] ), .B(\execute/alu/sll_175/ML_int[1][14] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][16] ) );
  MUX21 \execute/alu/sll_175/M1_1_12  ( .A(\execute/alu/sll_175/ML_int[1][12] ), .B(\execute/alu/sll_175/ML_int[1][10] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][12] ) );
  MUX21 \execute/alu/sll_175/M1_1_14  ( .A(\execute/alu/sll_175/ML_int[1][14] ), .B(\execute/alu/sll_175/ML_int[1][12] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][14] ) );
  MUX21 \execute/alu/sll_175/M1_0_22  ( .A(n1450), .B(n1449), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][22] ) );
  MUX21 \execute/alu/sll_175/M1_0_21  ( .A(n1449), .B(n1448), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][21] ) );
  MUX21 \execute/alu/sll_175/M1_0_30  ( .A(n1460), .B(n1458), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][30] ) );
  MUX21 \execute/alu/sll_175/M1_0_31  ( .A(n1461), .B(n1460), .S(
        \execute/alu/sll_175/temp_int_SH[0] ), .Q(
        \execute/alu/sll_175/ML_int[1][31] ) );
  MUX21 \execute/alu/sll_175/M1_1_31  ( .A(\execute/alu/sll_175/ML_int[1][31] ), .B(\execute/alu/sll_175/ML_int[1][29] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][31] ) );
  MUX21 \execute/alu/sll_175/M1_2_22  ( .A(\execute/alu/sll_175/ML_int[2][22] ), .B(\execute/alu/sll_175/ML_int[2][18] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][22] ) );
  MUX21 \execute/alu/sll_175/M1_2_18  ( .A(\execute/alu/sll_175/ML_int[2][18] ), .B(\execute/alu/sll_175/ML_int[2][14] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][18] ) );
  MUX21 \execute/alu/sll_175/M1_1_21  ( .A(\execute/alu/sll_175/ML_int[1][21] ), .B(\execute/alu/sll_175/ML_int[1][19] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][21] ) );
  MUX21 \execute/alu/sll_175/M1_2_4  ( .A(\execute/alu/sll_175/ML_int[2][4] ), 
        .B(\execute/alu/sll_175/ML_int[2][0] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][4] ) );
  MUX21 \execute/alu/sll_175/M1_2_20  ( .A(\execute/alu/sll_175/ML_int[2][20] ), .B(\execute/alu/sll_175/ML_int[2][16] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][20] ) );
  MUX21 \execute/alu/sll_175/M1_2_9  ( .A(\execute/alu/sll_175/ML_int[2][9] ), 
        .B(\execute/alu/sll_175/ML_int[2][5] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][9] ) );
  MUX21 \execute/alu/sll_175/M1_2_19  ( .A(\execute/alu/sll_175/ML_int[2][19] ), .B(\execute/alu/sll_175/ML_int[2][15] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][19] ) );
  MUX21 \execute/alu/sll_175/M1_2_11  ( .A(\execute/alu/sll_175/ML_int[2][11] ), .B(\execute/alu/sll_175/ML_int[2][7] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][11] ) );
  MUX21 \execute/alu/sll_175/M1_0_6  ( .A(n6193), .B(n1422), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][6] ) );
  MUX21 \execute/alu/sll_175/M1_0_24  ( .A(n1452), .B(n1451), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][24] ) );
  MUX21 \execute/alu/sll_175/M1_0_23  ( .A(n1451), .B(n1450), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][23] ) );
  MUX21 \execute/alu/sll_175/M1_0_29  ( .A(n1458), .B(n1457), .S(
        \execute/alu/sll_175/temp_int_SH[0] ), .Q(
        \execute/alu/sll_175/ML_int[1][29] ) );
  MUX21 \execute/alu/sll_175/M1_0_20  ( .A(n1448), .B(n1447), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][20] ) );
  MUX21 \execute/alu/sll_175/M1_0_17  ( .A(n1443), .B(n6222), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][17] ) );
  MUX21 \execute/alu/sll_175/M1_0_25  ( .A(n1453), .B(n1452), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][25] ) );
  MUX21 \execute/alu/sll_175/M1_0_8  ( .A(n1426), .B(n1425), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][8] ) );
  MUX21 \execute/alu/sll_175/M1_0_18  ( .A(n1445), .B(n1443), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][18] ) );
  MUX21 \execute/alu/sll_175/M1_0_27  ( .A(n1456), .B(n1454), .S(n6761), .Q(
        \execute/alu/sll_175/ML_int[1][27] ) );
  MUX21 \execute/alu/sll_175/M1_0_9  ( .A(n1427), .B(n1426), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][9] ) );
  MUX21 \execute/alu/sll_175/M1_0_28  ( .A(n1457), .B(n1456), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][28] ) );
  MUX21 \execute/alu/sll_175/M1_2_12  ( .A(\execute/alu/sll_175/ML_int[2][12] ), .B(\execute/alu/sll_175/ML_int[2][8] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][12] ) );
  MUX21 \execute/alu/sll_175/M1_0_26  ( .A(n1454), .B(n1453), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][26] ) );
  MUX21 \execute/alu/sll_175/M1_1_28  ( .A(\execute/alu/sll_175/ML_int[1][28] ), .B(\execute/alu/sll_175/ML_int[1][26] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][28] ) );
  MUX21 \execute/alu/sll_175/M1_2_28  ( .A(\execute/alu/sll_175/ML_int[2][28] ), .B(\execute/alu/sll_175/ML_int[2][24] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][28] ) );
  MUX21 \execute/alu/sll_175/M1_2_27  ( .A(\execute/alu/sll_175/ML_int[2][27] ), .B(\execute/alu/sll_175/ML_int[2][23] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][27] ) );
  MUX21 \execute/alu/sll_175/M1_1_29  ( .A(\execute/alu/sll_175/ML_int[1][29] ), .B(\execute/alu/sll_175/ML_int[1][27] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][29] ) );
  MUX21 \execute/alu/sll_175/M1_3_17  ( .A(\execute/alu/sll_175/ML_int[3][17] ), .B(\execute/alu/sll_175/ML_int[3][9] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][17] ) );
  MUX21 \execute/alu/sll_175/M1_1_30  ( .A(\execute/alu/sll_175/ML_int[1][30] ), .B(\execute/alu/sll_175/ML_int[1][28] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][30] ) );
  MUX21 \execute/alu/sll_175/M1_2_30  ( .A(\execute/alu/sll_175/ML_int[2][30] ), .B(\execute/alu/sll_175/ML_int[2][26] ), .S(n6758), .Q(
        \execute/alu/sll_175/ML_int[3][30] ) );
  MUX21 \execute/alu/sll_175/M1_4_30  ( .A(\execute/alu/sll_175/ML_int[4][30] ), .B(\execute/alu/sll_175/ML_int[4][14] ), .S(n6343), .Q(
        \execute/alu/sll_175/ML_int[5][30] ) );
  MUX21 \execute/alu/sll_175/M1_4_21  ( .A(\execute/alu/sll_175/ML_int[4][21] ), .B(n5809), .S(n6343), .Q(\execute/alu/sll_175/ML_int[5][21] ) );
  MUX21 \execute/alu/sll_175/M1_3_13  ( .A(\execute/alu/sll_175/ML_int[3][13] ), .B(\execute/alu/sll_175/ML_int[3][5] ), .S(n5819), .Q(
        \execute/alu/sll_175/ML_int[4][13] ) );
  MUX21 \execute/alu/sll_175/M1_1_25  ( .A(\execute/alu/sll_175/ML_int[1][25] ), .B(\execute/alu/sll_175/ML_int[1][23] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][25] ) );
  MUX21 \execute/alu/sll_175/M1_1_26  ( .A(\execute/alu/sll_175/ML_int[1][26] ), .B(\execute/alu/sll_175/ML_int[1][24] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][26] ) );
  MUX21 \execute/alu/sll_175/M1_1_27  ( .A(\execute/alu/sll_175/ML_int[1][27] ), .B(\execute/alu/sll_175/ML_int[1][25] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][27] ) );
  DF1 \memory/read_data_reg[1]  ( .D(ram_word[1]), .C(clk), .QN(n5642) );
  DF1 \memory/address_WB_reg[1]  ( .D(ram_adr[1]), .C(clk), .QN(n5643) );
  DF1 \instruction_decode/imm_reg[7]  ( .D(inst_out[7]), .C(clk), .Q(n6072) );
  DF3 \memory/address_WB_reg[21]  ( .D(ram_adr[21]), .C(clk), .QN(n5647) );
  DF3 \memory/address_WB_reg[10]  ( .D(ram_adr[10]), .C(clk), .QN(n5681) );
  DF3 \memory/address_WB_reg[20]  ( .D(ram_adr[20]), .C(clk), .QN(n5661) );
  MUX22 \execute/alu/sll_175/M1_2_21  ( .A(\execute/alu/sll_175/ML_int[2][21] ), .B(\execute/alu/sll_175/ML_int[2][17] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][21] ) );
  MUX22 \execute/alu/sll_175/M1_2_16  ( .A(\execute/alu/sll_175/ML_int[2][16] ), .B(\execute/alu/sll_175/ML_int[2][12] ), .S(n6757), .Q(
        \execute/alu/sll_175/ML_int[3][16] ) );
  DF1 \memory/address_WB_reg[16]  ( .D(ram_adr[16]), .C(clk), .QN(n5679) );
  DF1 \memory/address_WB_reg[17]  ( .D(ram_adr[17]), .C(clk), .QN(n5683) );
  MUX22 \execute/alu/sll_175/M1_1_15  ( .A(\execute/alu/sll_175/ML_int[1][15] ), .B(\execute/alu/sll_175/ML_int[1][13] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][15] ) );
  MUX22 \execute/alu/sll_175/M1_1_8  ( .A(\execute/alu/sll_175/ML_int[1][8] ), 
        .B(\execute/alu/sll_175/ML_int[1][6] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][8] ) );
  MUX22 \execute/alu/sll_175/M1_1_20  ( .A(\execute/alu/sll_175/ML_int[1][20] ), .B(\execute/alu/sll_175/ML_int[1][18] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][20] ) );
  MUX22 \execute/alu/sll_175/M1_1_10  ( .A(\execute/alu/sll_175/ML_int[1][10] ), .B(\execute/alu/sll_175/ML_int[1][8] ), .S(n5820), .Q(
        \execute/alu/sll_175/ML_int[2][10] ) );
  MUX22 \execute/alu/sll_175/M1_0_1  ( .A(n1415), .B(n1414), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][1] ) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[25][30]  ( .D(n6991), .E(
        n6808), .C(n1107), .RN(n6666), .QN(n4994) );
  MUX22 \execute/alu/sll_175/M1_0_7  ( .A(n1425), .B(n6193), .S(n6760), .Q(
        \execute/alu/sll_175/ML_int[1][7] ) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[25][21]  ( .D(
        write_data_reg[21]), .E(n6809), .C(n1107), .RN(n6665), .QN(n5164) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[25][27]  ( .D(n6985), .E(
        n6808), .C(n1107), .RN(n6665), .QN(n5334) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[15][29]  ( .D(n6989), .E(
        n6893), .C(n1107), .RN(n6676), .QN(n4840) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[25][29]  ( .D(n6989), .E(
        n6808), .C(n1107), .RN(n6666), .QN(n5044) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[27][27]  ( .D(n6985), .E(
        n6818), .C(n1107), .RN(n6662), .QN(n5174) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[24][30]  ( .D(n6991), .E(
        n6803), .C(n1107), .RN(n6618), .QN(n4995) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][29]  ( .D(n6989), .E(
        n6828), .C(n1107), .RN(n6659), .QN(n5040) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[27][28]  ( .D(n6987), .E(
        n6818), .C(n1107), .RN(n6662), .QN(n5118) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[11][30]  ( .D(n6991), .E(
        n6913), .C(n1107), .RN(n6683), .QN(n4954) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][2]  ( .D(n6934), .E(
        n6832), .C(n1107), .RN(n6656), .QN(n5194) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[15][2]  ( .D(
        write_data_reg[2]), .E(n6897), .C(n1107), .RN(n6673), .QN(n4868) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][12]  ( .D(
        write_data_reg[12]), .E(n6810), .C(n1107), .RN(n6664), .QN(n5210) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[25][1]  ( .D(n6932), .E(
        n6812), .C(n1107), .RN(n6663), .QN(n5302) );
  DFEC1 \instruction_decode/reg_MAPP/reg_file_reg[29][27]  ( .D(n6985), .E(
        n6828), .C(n1107), .RN(n6658), .QN(n5172) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[25][5]  ( .D(n6941), .E(
        n6811), .C(n1107), .RN(n6663), .QN(n5238) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[29][30]  ( .D(n6991), .E(
        n6828), .C(n1107), .RN(n6659), .QN(n4990) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[9][30]  ( .D(n6991), .E(
        n6903), .C(n1107), .RN(n6687), .QN(n4956) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[25][28]  ( .D(n6987), .E(
        n6808), .C(n1107), .RN(n6666), .QN(n5120) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[25][31]  ( .D(
        write_data_reg[31]), .E(n6808), .C(n1107), .RN(n6666), .QN(n5244) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[25][26]  ( .D(n6983), .E(
        n6808), .C(n1107), .RN(n6665), .QN(n5060) );
  DFEC3 \instruction_decode/reg_MAPP/reg_file_reg[27][2]  ( .D(n6934), .E(
        n6822), .C(n1107), .RN(n6659), .QN(n5196) );
  OAI221 U3767 ( .A(n4843), .B(n6587), .C(n4842), .D(n6583), .Q(n2996) );
  NOR42 U3768 ( .A(n2321), .B(n2322), .C(n2323), .D(n2324), .Q(n2320) );
  NAND43 U3769 ( .A(n1871), .B(n1872), .C(n1873), .D(n1874), .Q(n1870) );
  NOR41 U3770 ( .A(n3262), .B(n3263), .C(n3264), .D(n3265), .Q(n3261) );
  NOR41 U3771 ( .A(n2619), .B(n2620), .C(n2621), .D(n2622), .Q(n2613) );
  NOR41 U3772 ( .A(n3308), .B(n3309), .C(n3310), .D(n3311), .Q(n3302) );
  NOR42 U3773 ( .A(n3010), .B(n3011), .C(n3012), .D(n3013), .Q(n3009) );
  NOR42 U3774 ( .A(n2447), .B(n2448), .C(n2449), .D(n2450), .Q(n2446) );
  NOR41 U3775 ( .A(n2178), .B(n2179), .C(n2180), .D(n2181), .Q(n2172) );
  NOR41 U3776 ( .A(n2762), .B(n2763), .C(n2764), .D(n2765), .Q(n2756) );
  NOR41 U3777 ( .A(n2842), .B(n2843), .C(n2844), .D(n2845), .Q(n2841) );
  NOR41 U3778 ( .A(n2262), .B(n2263), .C(n2264), .D(n2265), .Q(n2256) );
  NOR42 U3779 ( .A(n3136), .B(n3137), .C(n3138), .D(n3139), .Q(n3135) );
  NOR42 U3780 ( .A(n3325), .B(n3326), .C(n3327), .D(n3328), .Q(n3324) );
  NOR42 U3781 ( .A(n2968), .B(n2969), .C(n2970), .D(n2971), .Q(n2967) );
  NOR42 U3782 ( .A(n3340), .B(n3341), .C(n3342), .D(n3343), .Q(n3339) );
  NOR42 U3783 ( .A(n2651), .B(n2652), .C(n2653), .D(n2654), .Q(n2650) );
  NOR42 U3784 ( .A(n2189), .B(n2190), .C(n2191), .D(n2192), .Q(n2188) );
  NOR42 U3785 ( .A(n2199), .B(n2200), .C(n2201), .D(n2202), .Q(n2193) );
  NOR42 U3786 ( .A(n1899), .B(n1900), .C(n1901), .D(n1902), .Q(n1893) );
  NOR41 U3787 ( .A(n2594), .B(n2595), .C(n2596), .D(n2597), .Q(n2593) );
  NOR42 U3788 ( .A(n2888), .B(n2889), .C(n2890), .D(n2891), .Q(n2882) );
  OAI221 U3789 ( .A(n4869), .B(n6551), .C(n4868), .D(n2009), .Q(n2223) );
  NOR41 U3790 ( .A(n2926), .B(n2927), .C(n2928), .D(n2929), .Q(n2925) );
  OAI221 U3791 ( .A(n5041), .B(n6578), .C(n5040), .D(n1928), .Q(n2928) );
  NOR23 U3792 ( .A(n2387), .B(n2386), .Q(n6108) );
  NOR42 U3793 ( .A(n2294), .B(n2295), .C(n2296), .D(n2297), .Q(n2293) );
  NOR42 U3794 ( .A(n2905), .B(n2906), .C(n2907), .D(n2908), .Q(n2904) );
  NOR23 U3795 ( .A(n2307), .B(n2306), .Q(n6118) );
  INV6 U3796 ( .A(rt[4]), .Q(n1490) );
  INV10 U3797 ( .A(n6486), .Q(n1143) );
  NOR41 U3798 ( .A(n2273), .B(n2274), .C(n2275), .D(n2276), .Q(n2272) );
  INV3 U3799 ( .A(n6334), .Q(n5814) );
  INV3 U3800 ( .A(n5814), .Q(n5815) );
  INV3 U3801 ( .A(n5814), .Q(n5816) );
  NAND24 U3802 ( .A(n1320), .B(n4248), .Q(n3589) );
  AOI212 U3803 ( .A(n3690), .B(n3936), .C(n4244), .Q(n4246) );
  NOR41 U3804 ( .A(n4308), .B(n4309), .C(n4310), .D(n1388), .Q(n4307) );
  INV6 U3805 ( .A(n4444), .Q(n1449) );
  NOR42 U3806 ( .A(n2279), .B(n2280), .C(n2281), .D(n2282), .Q(n2278) );
  AOI222 U3807 ( .A(ram_adr[9]), .B(n6337), .C(n6339), .D(data_1[9]), .Q(n4534) );
  NOR33 U3808 ( .A(n6201), .B(n4048), .C(n4049), .Q(n4046) );
  OAI222 U3809 ( .A(n3542), .B(n3515), .C(n3477), .D(n3476), .Q(n4243) );
  NAND28 U3810 ( .A(n6194), .B(n6195), .Q(n3476) );
  INV6 U3811 ( .A(n4139), .Q(n1369) );
  INV6 U3812 ( .A(n6264), .Q(n1311) );
  AOI210 U3813 ( .A(n6512), .B(n3592), .C(n3594), .Q(n3578) );
  AOI220 U3814 ( .A(n1470), .B(n1338), .C(n6515), .D(n3592), .Q(n3583) );
  OAI2110 U3815 ( .A(n3592), .B(n6514), .C(n3593), .D(n6352), .Q(n3585) );
  NAND20 U3816 ( .A(n6516), .B(n3592), .Q(n3593) );
  CLKBU4 U3817 ( .A(\execute/alu/sll_175/temp_int_SH[0] ), .Q(n6761) );
  CLKBU4 U3818 ( .A(\execute/alu/sll_175/temp_int_SH[0] ), .Q(n6760) );
  NAND21 U3819 ( .A(n4020), .B(n1383), .Q(n4003) );
  XNR22 U3820 ( .A(n4018), .B(n6350), .Q(n4020) );
  NOR21 U3821 ( .A(n3806), .B(n1404), .Q(n3739) );
  BUF6 U3822 ( .A(n3683), .Q(n5817) );
  CLKIN6 U3823 ( .A(\execute/op_21 [12]), .Q(n1433) );
  NAND22 U3824 ( .A(n6222), .B(n6321), .Q(n6224) );
  INV6 U3825 ( .A(n4039), .Q(n6222) );
  INV3 U3826 ( .A(\execute/alu/sll_175/temp_int_SH[3] ), .Q(n5818) );
  INV3 U3827 ( .A(n5818), .Q(n5819) );
  OAI210 U3828 ( .A(n4458), .B(n1338), .C(n4401), .Q(
        \execute/alu/sll_175/temp_int_SH[3] ) );
  OAI212 U3829 ( .A(n4056), .B(n4048), .C(n4057), .Q(n4045) );
  NOR22 U3830 ( .A(n4111), .B(n4110), .Q(n4048) );
  NOR41 U3831 ( .A(n3277), .B(n3278), .C(n3279), .D(n3280), .Q(n3276) );
  NAND20 U3832 ( .A(n4054), .B(n4053), .Q(n3561) );
  NOR22 U3833 ( .A(n1975), .B(n1982), .Q(\instruction_decode/old_ex [1]) );
  AOI220 U3834 ( .A(n1470), .B(n1320), .C(n6515), .D(n5817), .Q(n3685) );
  NOR20 U3835 ( .A(n5817), .B(n3404), .Q(n3684) );
  NAND20 U3836 ( .A(n5817), .B(n3592), .Q(n3604) );
  INV10 U3837 ( .A(n5817), .Q(n1320) );
  OAI210 U3838 ( .A(n5716), .B(n1969), .C(n1970), .Q(
        \instruction_decode/old_m [3]) );
  NAND33 U3839 ( .A(n1773), .B(n5945), .C(n5717), .Q(n1970) );
  CLKBU15 U3840 ( .A(\execute/n434 ), .Q(n5829) );
  OAI2112 U3841 ( .A(n3850), .B(n3870), .C(n4303), .D(n4304), .Q(n4301) );
  NAND26 U3842 ( .A(n6489), .B(\execute/op_21 [22]), .Q(n3870) );
  BUF6 U3843 ( .A(\execute/alu/sll_175/temp_int_SH[1] ), .Q(n5820) );
  XNR21 U3844 ( .A(n1472), .B(n3930), .Q(n3691) );
  CLKIN4 U3845 ( .A(n3930), .Q(n1415) );
  NOR22 U3846 ( .A(n3910), .B(n1393), .Q(n3872) );
  BUF2 U3847 ( .A(n4134), .Q(n5821) );
  OAI210 U3848 ( .A(n3938), .B(n6341), .C(n6321), .Q(n3937) );
  OAI210 U3849 ( .A(n3938), .B(n6341), .C(n3936), .Q(n4380) );
  NAND26 U3850 ( .A(n3938), .B(n6341), .Q(n3936) );
  XNR22 U3851 ( .A(n6350), .B(n1414), .Q(n3938) );
  NAND26 U3852 ( .A(n1372), .B(n4130), .Q(n4058) );
  XNR22 U3853 ( .A(n1472), .B(n6346), .Q(n4130) );
  INV3 U3854 ( .A(n4549), .Q(n5822) );
  CLKIN6 U3855 ( .A(n5822), .Q(n5823) );
  NOR23 U3856 ( .A(n6235), .B(n4394), .Q(n6236) );
  NAND43 U3857 ( .A(n4469), .B(n4470), .C(n4471), .D(n4472), .Q(n4394) );
  AOI220 U3858 ( .A(n5944), .B(n6490), .C(\execute/op_21 [6]), .D(n6489), .Q(
        n5824) );
  AOI222 U3859 ( .A(n5944), .B(n6490), .C(\execute/op_21 [6]), .D(n6489), .Q(
        n3508) );
  BUF15 U3860 ( .A(n3508), .Q(n6348) );
  INV15 U3861 ( .A(n6348), .Q(n6193) );
  NOR41 U3862 ( .A(n1875), .B(n1876), .C(n1877), .D(n1878), .Q(n1874) );
  XOR21 U3863 ( .A(\instruction_decode/old_data_2 [13]), .B(
        \instruction_decode/reg_MAPP/n3641 ), .Q(n1876) );
  INV3 U3864 ( .A(n4291), .Q(n6335) );
  NOR40 U3865 ( .A(n3203), .B(n3204), .C(n3205), .D(n3206), .Q(n3197) );
  NOR40 U3866 ( .A(n2493), .B(n2494), .C(n2495), .D(n2496), .Q(n2487) );
  INV3 U3867 ( .A(n3740), .Q(n1407) );
  NOR21 U3868 ( .A(n3662), .B(n3657), .Q(n3631) );
  NOR21 U3869 ( .A(n3185), .B(n3184), .Q(n6152) );
  NOR21 U3870 ( .A(n3227), .B(n3226), .Q(n6154) );
  NOR21 U3871 ( .A(n3269), .B(n3268), .Q(n6179) );
  NOR21 U3872 ( .A(n2744), .B(n2743), .Q(n6172) );
  NOR21 U3873 ( .A(n2601), .B(n2600), .Q(n6150) );
  NOR21 U3874 ( .A(n2019), .B(n2018), .Q(n6174) );
  NOR21 U3875 ( .A(n2139), .B(n2138), .Q(n6185) );
  NOR21 U3876 ( .A(n2685), .B(n2684), .Q(n6160) );
  INV6 U3877 ( .A(n6283), .Q(n6284) );
  INV6 U3878 ( .A(n3592), .Q(n1338) );
  CLKIN12 U3879 ( .A(n6338), .Q(n6340) );
  CLKIN4 U3880 ( .A(n6335), .Q(n6336) );
  NOR40 U3881 ( .A(n1921), .B(n1922), .C(n1923), .D(n1924), .Q(n1920) );
  INV3 U3882 ( .A(n6130), .Q(n6131) );
  NOR40 U3883 ( .A(n2510), .B(n2511), .C(n2512), .D(n2513), .Q(n2509) );
  INV3 U3884 ( .A(n6134), .Q(n6135) );
  NOR40 U3885 ( .A(n2573), .B(n2574), .C(n2575), .D(n2576), .Q(n2572) );
  NOR40 U3886 ( .A(n2069), .B(n2070), .C(n2071), .D(n2072), .Q(n2068) );
  NOR40 U3887 ( .A(n2153), .B(n2154), .C(n2155), .D(n2156), .Q(n2152) );
  INV3 U3888 ( .A(n6116), .Q(n6117) );
  INV3 U3889 ( .A(n6239), .Q(n6240) );
  NOR21 U3890 ( .A(n6188), .B(n3049), .Q(n3045) );
  NOR21 U3891 ( .A(n6184), .B(n3112), .Q(n3108) );
  NOR21 U3892 ( .A(n6127), .B(n3154), .Q(n3150) );
  NOR21 U3893 ( .A(n6137), .B(n3175), .Q(n3171) );
  NOR41 U3894 ( .A(n3193), .B(n3194), .C(n3195), .D(n3196), .Q(n3192) );
  NOR21 U3895 ( .A(n6139), .B(n3217), .Q(n3213) );
  NOR21 U3896 ( .A(n6165), .B(n3259), .Q(n3255) );
  NOR41 U3897 ( .A(n3319), .B(n3320), .C(n3321), .D(n3322), .Q(n3318) );
  NOR41 U3898 ( .A(n2710), .B(n2711), .C(n2712), .D(n2713), .Q(n2709) );
  NOR21 U3899 ( .A(n6157), .B(n2734), .Q(n2730) );
  NOR21 U3900 ( .A(n6192), .B(n2839), .Q(n2835) );
  NOR41 U3901 ( .A(n2336), .B(n2337), .C(n2338), .D(n2339), .Q(n2335) );
  NOR41 U3902 ( .A(n2357), .B(n2358), .C(n2359), .D(n2360), .Q(n2356) );
  NOR21 U3903 ( .A(n6182), .B(n2465), .Q(n2461) );
  NOR41 U3904 ( .A(n2483), .B(n2484), .C(n2485), .D(n2486), .Q(n2482) );
  NOR21 U3905 ( .A(n6133), .B(n2591), .Q(n2587) );
  NOR21 U3906 ( .A(n6159), .B(n2001), .Q(n1997) );
  NOR41 U3907 ( .A(n2042), .B(n2043), .C(n2044), .D(n2045), .Q(n2041) );
  NOR21 U3908 ( .A(n6167), .B(n2129), .Q(n2125) );
  NOR21 U3909 ( .A(n6141), .B(n2675), .Q(n2671) );
  AOI2111 U3910 ( .A(n3477), .B(n6348), .C(n4324), .D(n4325), .Q(n4322) );
  NAND23 U3911 ( .A(n1370), .B(n4165), .Q(n4139) );
  NAND42 U3912 ( .A(n4552), .B(n1728), .C(n4553), .D(n4554), .Q(n4543) );
  INV3 U3913 ( .A(n6245), .Q(n4417) );
  NAND22 U3914 ( .A(n5733), .B(n6217), .Q(n6216) );
  INV3 U3915 ( .A(n6231), .Q(n4409) );
  NAND22 U3916 ( .A(n6246), .B(n6232), .Q(n6231) );
  NAND22 U3917 ( .A(n6267), .B(n4479), .Q(n4541) );
  NOR21 U3918 ( .A(n4165), .B(n1370), .Q(n4059) );
  INV3 U3919 ( .A(n4058), .Q(n1371) );
  INV3 U3920 ( .A(n6218), .Q(n6219) );
  OAI311 U3921 ( .A(n3633), .B(n3631), .C(n1380), .D(n3635), .Q(n3629) );
  AOI311 U3922 ( .A(n3639), .B(n3640), .C(n3641), .D(n3642), .Q(n3638) );
  INV3 U3923 ( .A(n6216), .Q(n1986) );
  NOR21 U3924 ( .A(n1936), .B(n1934), .Q(n6130) );
  INV3 U3925 ( .A(n6096), .Q(n6097) );
  NOR21 U3926 ( .A(n3290), .B(n3289), .Q(n6096) );
  INV3 U3927 ( .A(n6118), .Q(n6119) );
  NOR21 U3928 ( .A(n2517), .B(n2516), .Q(n6134) );
  NOR21 U3929 ( .A(n2160), .B(n2159), .Q(n6116) );
  NAND31 U3930 ( .A(reg_write), .B(n5943), .C(write_register[3]), .Q(n1955) );
  NAND31 U3931 ( .A(write_register[4]), .B(reg_write), .C(write_register[3]), 
        .Q(n1965) );
  NAND31 U3932 ( .A(n6069), .B(n5943), .C(reg_write), .Q(n1966) );
  NAND31 U3933 ( .A(reg_write), .B(n6069), .C(write_register[4]), .Q(n1964) );
  INV3 U3934 ( .A(n6220), .Q(n6221) );
  AOI221 U3935 ( .A(ram_adr[1]), .B(n6337), .C(n6340), .D(data_1[1]), .Q(n4467) );
  INV8 U3936 ( .A(n6347), .Q(n1420) );
  INV3 U3937 ( .A(n3528), .Q(n1351) );
  INV3 U3938 ( .A(n3542), .Q(n1356) );
  INV6 U3939 ( .A(n3465), .Q(n1425) );
  NAND22 U3940 ( .A(n3476), .B(n3477), .Q(n3475) );
  NAND22 U3941 ( .A(n1472), .B(n5824), .Q(n6194) );
  NAND24 U3942 ( .A(n6351), .B(n6193), .Q(n6195) );
  OAI2111 U3943 ( .A(n6940), .B(n6505), .C(n4459), .D(n4460), .Q(n3564) );
  NAND26 U3944 ( .A(n6177), .B(n6178), .Q(n4171) );
  NAND22 U3945 ( .A(n6176), .B(n6344), .Q(n6178) );
  NAND23 U3946 ( .A(n1472), .B(n1430), .Q(n6177) );
  INV3 U3947 ( .A(n4175), .Q(n1429) );
  INV3 U3948 ( .A(n4256), .Q(n1258) );
  NOR22 U3949 ( .A(n3976), .B(n1381), .Q(n4002) );
  NOR21 U3950 ( .A(n1446), .B(n3998), .Q(n3974) );
  NAND23 U3951 ( .A(n1338), .B(n1320), .Q(n3601) );
  NAND22 U3952 ( .A(n6207), .B(n6208), .Q(n3875) );
  NAND22 U3953 ( .A(n4444), .B(n6350), .Q(n6208) );
  NAND23 U3954 ( .A(n3875), .B(n1395), .Q(n3874) );
  BUF2 U3955 ( .A(n1472), .Q(n6322) );
  XNR21 U3956 ( .A(n3843), .B(n6350), .Q(n3827) );
  INV6 U3957 ( .A(n6198), .Q(n6199) );
  NAND22 U3958 ( .A(n3737), .B(n1408), .Q(n3740) );
  INV3 U3959 ( .A(n6335), .Q(n6337) );
  INV3 U3960 ( .A(n3611), .Q(n1293) );
  INV3 U3961 ( .A(n3610), .Q(n1289) );
  INV3 U3962 ( .A(n6338), .Q(n6339) );
  INV3 U3963 ( .A(n4572), .Q(n1728) );
  OAI311 U3964 ( .A(write_register_ex[0]), .B(write_register_ex[1]), .C(n6225), 
        .D(wb_MEM[1]), .Q(n4572) );
  NAND33 U3965 ( .A(n6226), .B(n6268), .C(n6227), .Q(n6225) );
  XNR21 U3966 ( .A(write_register_ex[4]), .B(n1490), .Q(n4569) );
  NAND23 U3967 ( .A(n4566), .B(n4567), .Q(n6144) );
  OAI311 U3968 ( .A(n1960), .B(write_register[4]), .C(write_register[3]), .D(
        reg_write), .Q(n4549) );
  NOR40 U3969 ( .A(n2930), .B(n2931), .C(n2932), .D(n2933), .Q(n2924) );
  NOR40 U3970 ( .A(n3052), .B(n3053), .C(n3054), .D(n3055), .Q(n3051) );
  NOR40 U3971 ( .A(n3056), .B(n3057), .C(n3058), .D(n3059), .Q(n3050) );
  NOR40 U3972 ( .A(n3115), .B(n3116), .C(n3117), .D(n3118), .Q(n3114) );
  NOR40 U3973 ( .A(n3119), .B(n3120), .C(n3121), .D(n3122), .Q(n3113) );
  NOR40 U3974 ( .A(n3157), .B(n3158), .C(n3159), .D(n3160), .Q(n3156) );
  NOR40 U3975 ( .A(n3178), .B(n3179), .C(n3180), .D(n3181), .Q(n3177) );
  INV3 U3976 ( .A(n6152), .Q(n6153) );
  NOR40 U3977 ( .A(n3220), .B(n3221), .C(n3222), .D(n3223), .Q(n3219) );
  INV3 U3978 ( .A(n6154), .Q(n6155) );
  INV3 U3979 ( .A(n6179), .Q(n6180) );
  NOR40 U3980 ( .A(n2737), .B(n2738), .C(n2739), .D(n2740), .Q(n2736) );
  INV3 U3981 ( .A(n6172), .Q(n6173) );
  NOR40 U3982 ( .A(n2846), .B(n2847), .C(n2848), .D(n2849), .Q(n2840) );
  INV3 U3983 ( .A(n6108), .Q(n6109) );
  NOR40 U3984 ( .A(n2468), .B(n2469), .C(n2470), .D(n2471), .Q(n2467) );
  INV3 U3985 ( .A(n6150), .Q(n6151) );
  INV3 U3986 ( .A(n6174), .Q(n6175) );
  NOR40 U3987 ( .A(n2004), .B(n2005), .C(n2006), .D(n2007), .Q(n2003) );
  INV3 U3988 ( .A(n6185), .Q(n6186) );
  NOR40 U3989 ( .A(n2132), .B(n2133), .C(n2134), .D(n2135), .Q(n2131) );
  NOR40 U3990 ( .A(n2220), .B(n2221), .C(n2222), .D(n2223), .Q(n2214) );
  NOR40 U3991 ( .A(n2216), .B(n2217), .C(n2218), .D(n2219), .Q(n2215) );
  NOR40 U3992 ( .A(n2678), .B(n2679), .C(n2680), .D(n2681), .Q(n2677) );
  INV3 U3993 ( .A(n6160), .Q(n6161) );
  INV6 U3994 ( .A(n5825), .Q(n5826) );
  INV3 U3995 ( .A(n6488), .Q(n5825) );
  INV3 U3996 ( .A(n6296), .Q(n6301) );
  AOI221 U3997 ( .A(ram_adr[2]), .B(n6336), .C(n6340), .D(data_1[2]), .Q(n4465) );
  NAND22 U3998 ( .A(n4533), .B(n4534), .Q(n3398) );
  AOI221 U3999 ( .A(n6503), .B(write_data_reg[9]), .C(pc_ex[9]), .D(n6324), 
        .Q(n4533) );
  AOI221 U4000 ( .A(n3859), .B(n4066), .C(\execute/alu/sll_175/ML_int[5][16] ), 
        .D(n1353), .Q(n4030) );
  BUF6 U4001 ( .A(\execute/n433 ), .Q(n5830) );
  INV3 U4002 ( .A(n1991), .Q(n1413) );
  NOR22 U4003 ( .A(n1983), .B(n1967), .Q(n1866) );
  NAND31 U4004 ( .A(n1985), .B(n5868), .C(n6085), .Q(n1973) );
  NOR21 U4005 ( .A(n6113), .B(n1918), .Q(n1914) );
  NOR40 U4006 ( .A(n2752), .B(n2753), .C(n2754), .D(n2755), .Q(n2751) );
  NOR41 U4007 ( .A(n2168), .B(n2169), .C(n2170), .D(n2171), .Q(n2167) );
  NOR41 U4008 ( .A(n2252), .B(n2253), .C(n2254), .D(n2255), .Q(n2251) );
  NOR41 U4009 ( .A(n2399), .B(n2400), .C(n2401), .D(n2402), .Q(n2398) );
  NOR41 U4010 ( .A(n2420), .B(n2421), .C(n2422), .D(n2423), .Q(n2419) );
  NOR21 U4011 ( .A(n6115), .B(n2507), .Q(n2503) );
  NOR40 U4012 ( .A(n2546), .B(n2547), .C(n2548), .D(n2549), .Q(n2545) );
  NOR21 U4013 ( .A(n6121), .B(n2570), .Q(n2566) );
  NOR21 U4014 ( .A(n6125), .B(n2066), .Q(n2062) );
  NOR21 U4015 ( .A(n6099), .B(n2150), .Q(n2146) );
  NOR40 U4016 ( .A(n4277), .B(n4278), .C(n1354), .D(n4279), .Q(n4276) );
  AOI221 U4017 ( .A(n6333), .B(data_2[16]), .C(n5815), .D(ram_adr[16]), .Q(
        n4451) );
  AOI221 U4018 ( .A(n6333), .B(data_2[13]), .C(n5815), .D(ram_adr[13]), .Q(
        n4454) );
  AOI221 U4019 ( .A(n6330), .B(data_2[10]), .C(n5815), .D(ram_adr[10]), .Q(
        n4457) );
  NAND33 U4020 ( .A(n4421), .B(n6267), .C(n4422), .Q(n5813) );
  NAND23 U4021 ( .A(n2856), .B(n6163), .Q(\instruction_decode/old_data_1 [31])
         );
  NAND42 U4022 ( .A(n2916), .B(n2917), .C(n2918), .D(n2919), .Q(
        \instruction_decode/old_data_1 [29]) );
  NAND22 U4023 ( .A(n3003), .B(n6143), .Q(\instruction_decode/old_data_1 [25])
         );
  NAND42 U4024 ( .A(n3042), .B(n3043), .C(n3044), .D(n3045), .Q(
        \instruction_decode/old_data_1 [23]) );
  NAND42 U4025 ( .A(n3105), .B(n3106), .C(n3107), .D(n3108), .Q(
        \instruction_decode/old_data_1 [20]) );
  NAND42 U4026 ( .A(n3147), .B(n3148), .C(n3149), .D(n3150), .Q(
        \instruction_decode/old_data_1 [19]) );
  NAND42 U4027 ( .A(n3168), .B(n3169), .C(n3170), .D(n3171), .Q(
        \instruction_decode/old_data_1 [18]) );
  NAND42 U4028 ( .A(n3189), .B(n3190), .C(n3191), .D(n3192), .Q(
        \instruction_decode/old_data_1 [17]) );
  NAND42 U4029 ( .A(n3210), .B(n3211), .C(n3212), .D(n3213), .Q(
        \instruction_decode/old_data_1 [16]) );
  NAND42 U4030 ( .A(n3252), .B(n3253), .C(n3254), .D(n3255), .Q(
        \instruction_decode/old_data_1 [14]) );
  NAND42 U4031 ( .A(n3315), .B(n3316), .C(n3317), .D(n3318), .Q(
        \instruction_decode/old_data_1 [10]) );
  NAND42 U4032 ( .A(n2706), .B(n2707), .C(n2708), .D(n2709), .Q(
        \instruction_decode/old_data_1 [9]) );
  NAND42 U4033 ( .A(n2727), .B(n2728), .C(n2729), .D(n2730), .Q(
        \instruction_decode/old_data_1 [8]) );
  NAND42 U4034 ( .A(n2832), .B(n2833), .C(n2834), .D(n2835), .Q(
        \instruction_decode/old_data_1 [3]) );
  NAND42 U4035 ( .A(n2311), .B(n2312), .C(n2313), .D(n2314), .Q(
        \instruction_decode/old_data_2 [25]) );
  NAND42 U4036 ( .A(n2332), .B(n2333), .C(n2334), .D(n2335), .Q(
        \instruction_decode/old_data_2 [24]) );
  NAND42 U4037 ( .A(n2353), .B(n2354), .C(n2355), .D(n2356), .Q(
        \instruction_decode/old_data_2 [23]) );
  NAND22 U4038 ( .A(n2377), .B(n6101), .Q(\instruction_decode/old_data_2 [22])
         );
  NAND42 U4039 ( .A(n2458), .B(n2459), .C(n2460), .D(n2461), .Q(
        \instruction_decode/old_data_2 [19]) );
  NAND42 U4040 ( .A(n2479), .B(n2480), .C(n2481), .D(n2482), .Q(
        \instruction_decode/old_data_2 [18]) );
  NAND42 U4041 ( .A(n2584), .B(n2585), .C(n2586), .D(n2587), .Q(
        \instruction_decode/old_data_2 [13]) );
  NAND42 U4042 ( .A(n1994), .B(n1995), .C(n1996), .D(n1997), .Q(
        \instruction_decode/old_data_2 [9]) );
  NAND42 U4043 ( .A(n2038), .B(n2039), .C(n2040), .D(n2041), .Q(
        \instruction_decode/old_data_2 [8]) );
  NAND42 U4044 ( .A(n2101), .B(n2102), .C(n2103), .D(n2104), .Q(
        \instruction_decode/old_data_2 [5]) );
  NAND42 U4045 ( .A(n2122), .B(n2123), .C(n2124), .D(n2125), .Q(
        \instruction_decode/old_data_2 [4]) );
  NAND42 U4046 ( .A(n2206), .B(n2207), .C(n2208), .D(n2209), .Q(
        \instruction_decode/old_data_2 [2]) );
  NAND42 U4047 ( .A(n2437), .B(n2438), .C(n2439), .D(n2440), .Q(
        \instruction_decode/old_data_2 [1]) );
  NAND42 U4048 ( .A(n2668), .B(n2669), .C(n2670), .D(n2671), .Q(
        \instruction_decode/old_data_2 [0]) );
  NOR42 U4049 ( .A(n3346), .B(n3347), .C(n3348), .D(n3349), .Q(n3345) );
  INV3 U4050 ( .A(\execute/op_21 [11]), .Q(n1431) );
  OAI221 U4051 ( .A(n6928), .B(n5690), .C(n6923), .D(n5691), .Q(
        write_data_reg[30]) );
  INV3 U4052 ( .A(\execute/op_21 [4]), .Q(n1421) );
  NOR42 U4053 ( .A(n3073), .B(n3074), .C(n3075), .D(n3076), .Q(n3072) );
  NOR42 U4054 ( .A(n3094), .B(n3095), .C(n3096), .D(n3097), .Q(n3093) );
  NAND26 U4055 ( .A(n1148), .B(n5717), .Q(n1974) );
  NAND23 U4056 ( .A(n1148), .B(n1980), .Q(n1979) );
  INV12 U4057 ( .A(n3681), .Q(n1416) );
  CLKBU15 U4058 ( .A(\execute/n431 ), .Q(n6345) );
  OAI220 U4059 ( .A(n4236), .B(n3398), .C(n4337), .D(n4325), .Q(n4321) );
  NAND20 U4060 ( .A(n3398), .B(n4236), .Q(n3421) );
  CLKIN1 U4061 ( .A(n4236), .Q(n1427) );
  INV3 U4062 ( .A(n6925), .Q(n5827) );
  INV3 U4063 ( .A(n5827), .Q(n5828) );
  INV0 U4064 ( .A(n6068), .Q(n6925) );
  INV3 U4065 ( .A(n3632), .Q(n6213) );
  BUF15 U4066 ( .A(n6326), .Q(n5831) );
  BUF15 U4067 ( .A(n6326), .Q(n5832) );
  CLKIN6 U4068 ( .A(n6325), .Q(n6326) );
  BUF12 U4069 ( .A(n3627), .Q(n6350) );
  NAND22 U4070 ( .A(n6516), .B(n6321), .Q(n3438) );
  OAI222 U4071 ( .A(n6926), .B(n5640), .C(n5828), .D(n5641), .Q(
        write_data_reg[2]) );
  CLKIN2 U4072 ( .A(n6935), .Q(n6934) );
  OAI222 U4073 ( .A(n6926), .B(n5642), .C(n5828), .D(n5643), .Q(
        write_data_reg[1]) );
  CLKIN2 U4074 ( .A(n6933), .Q(n6932) );
  OAI222 U4075 ( .A(n6926), .B(n5644), .C(n5828), .D(n5645), .Q(
        write_data_reg[4]) );
  CLKIN2 U4076 ( .A(n6940), .Q(n6939) );
  OAI222 U4077 ( .A(n6928), .B(n5658), .C(n6923), .D(n5659), .Q(
        write_data_reg[0]) );
  CLKIN2 U4078 ( .A(n6931), .Q(n6930) );
  INV3 U4079 ( .A(write_data_reg[29]), .Q(n6990) );
  INV3 U4080 ( .A(write_data_reg[30]), .Q(n6992) );
  INV3 U4081 ( .A(write_data_reg[28]), .Q(n6988) );
  INV3 U4082 ( .A(write_data_reg[25]), .Q(n6982) );
  NOR21 U4083 ( .A(n6265), .B(n1468), .Q(n6334) );
  INV12 U4084 ( .A(n6350), .Q(n1472) );
  INV3 U4085 ( .A(n6236), .Q(n3596) );
  INV3 U4086 ( .A(n4288), .Q(n1468) );
  CLKIN2 U4087 ( .A(n6286), .Q(n6307) );
  INV3 U4088 ( .A(write_data_reg[9]), .Q(n6950) );
  INV2 U4089 ( .A(n6327), .Q(n6328) );
  CLKIN3 U4090 ( .A(n6328), .Q(n6329) );
  OAI210 U4091 ( .A(n4458), .B(n1320), .C(n4401), .Q(
        \execute/alu/sll_175/temp_int_SH[2] ) );
  INV3 U4092 ( .A(\execute/alu/sll_175/temp_int_SH[2] ), .Q(n6759) );
  INV6 U4093 ( .A(n4427), .Q(n6331) );
  CLKIN6 U4094 ( .A(n6331), .Q(n6332) );
  CLKIN1 U4095 ( .A(n1486), .Q(n6265) );
  INV3 U4096 ( .A(n4425), .Q(n6325) );
  INV8 U4097 ( .A(n6344), .Q(n1430) );
  BUF8 U4098 ( .A(\execute/n430 ), .Q(n6344) );
  BUF12 U4099 ( .A(\execute/n453 ), .Q(n6347) );
  INV3 U4100 ( .A(n6281), .Q(n6308) );
  INV6 U4101 ( .A(n4424), .Q(n1484) );
  NAND23 U4102 ( .A(n4563), .B(n6107), .Q(n4424) );
  INV3 U4103 ( .A(n6942), .Q(n6941) );
  INV6 U4104 ( .A(n6964), .Q(n6963) );
  INV6 U4105 ( .A(n6954), .Q(n6953) );
  INV3 U4106 ( .A(n6976), .Q(n6975) );
  INV3 U4107 ( .A(n6944), .Q(n6943) );
  INV6 U4108 ( .A(n6962), .Q(n6961) );
  INV6 U4109 ( .A(n6958), .Q(n6957) );
  INV3 U4110 ( .A(n6759), .Q(n6757) );
  INV3 U4111 ( .A(n5819), .Q(n6756) );
  INV6 U4112 ( .A(n6345), .Q(n6210) );
  INV3 U4113 ( .A(n6253), .Q(n4039) );
  NAND31 U4114 ( .A(n6351), .B(n4343), .C(n4064), .Q(n3404) );
  OAI222 U4115 ( .A(n4921), .B(n6588), .C(n4920), .D(n1926), .Q(n2908) );
  NOR42 U4116 ( .A(n1879), .B(n1880), .C(n1881), .D(n1882), .Q(n1873) );
  NOR41 U4117 ( .A(n2962), .B(n2963), .C(n2964), .D(n2965), .Q(n2961) );
  NAND42 U4118 ( .A(n2269), .B(n2270), .C(n2271), .D(n2272), .Q(
        \instruction_decode/old_data_2 [27]) );
  NOR41 U4119 ( .A(n2237), .B(n2238), .C(n2239), .D(n2240), .Q(n2236) );
  NOR41 U4120 ( .A(n2231), .B(n2232), .C(n2233), .D(n2234), .Q(n2230) );
  NAND31 U4121 ( .A(n3128), .B(n3126), .C(n3127), .Q(n6092) );
  NAND22 U4122 ( .A(n3129), .B(n6093), .Q(\instruction_decode/old_data_1 [1])
         );
  INV3 U4123 ( .A(n6092), .Q(n6093) );
  NOR41 U4124 ( .A(n3130), .B(n3131), .C(n3132), .D(n3133), .Q(n3129) );
  OAI222 U4125 ( .A(n5163), .B(n6532), .C(n5162), .D(n6527), .Q(n2406) );
  NAND31 U4126 ( .A(n2876), .B(n2874), .C(n2875), .Q(n6094) );
  NAND22 U4127 ( .A(n2877), .B(n6095), .Q(\instruction_decode/old_data_1 [30])
         );
  INV3 U4128 ( .A(n6094), .Q(n6095) );
  NOR41 U4129 ( .A(n2878), .B(n2879), .C(n2880), .D(n2881), .Q(n2877) );
  OAI222 U4130 ( .A(n5009), .B(n6531), .C(n5008), .D(n2013), .Q(n2410) );
  NOR22 U4131 ( .A(n2244), .B(n2243), .Q(n6128) );
  INV4 U4132 ( .A(n6283), .Q(n6278) );
  INV10 U4133 ( .A(n6310), .Q(n6283) );
  BUF15 U4134 ( .A(n1777), .Q(n6486) );
  NAND28 U4135 ( .A(n6284), .B(n6270), .Q(n1777) );
  NOR42 U4136 ( .A(n1895), .B(n1896), .C(n1897), .D(n1898), .Q(n1894) );
  NOR22 U4137 ( .A(n6309), .B(n1125), .Q(n5751) );
  CLKIN2 U4138 ( .A(n6308), .Q(n6309) );
  OAI211 U4139 ( .A(n5826), .B(n1155), .C(n1832), .Q(n5795) );
  AOI221 U4140 ( .A(n1833), .B(n6313), .C(n1142), .D(inst_out[9]), .Q(n1832)
         );
  INV4 U4141 ( .A(n6278), .Q(n6313) );
  INV2 U4142 ( .A(n6310), .Q(n6311) );
  INV3 U4143 ( .A(n6278), .Q(n6314) );
  OAI222 U4144 ( .A(n5323), .B(n6522), .C(n5322), .D(n6519), .Q(n2409) );
  OAI211 U4145 ( .A(n5826), .B(n1159), .C(n1782), .Q(n5776) );
  OAI211 U4146 ( .A(n6487), .B(n1158), .C(n1797), .Q(n5782) );
  OAI211 U4147 ( .A(n6487), .B(n1154), .C(n1778), .Q(n5775) );
  OAI211 U4148 ( .A(n6487), .B(n5706), .C(n1785), .Q(n5777) );
  OAI211 U4149 ( .A(n6487), .B(n5704), .C(n1791), .Q(n5779) );
  OAI211 U4150 ( .A(n6487), .B(n5705), .C(n1823), .Q(n5792) );
  CLKIN6 U4151 ( .A(n6270), .Q(n1142) );
  NOR42 U4152 ( .A(n1371), .B(n4062), .C(n1369), .D(n4063), .Q(n4060) );
  NAND26 U4153 ( .A(n1987), .B(n6242), .Q(n1768) );
  INV2 U4154 ( .A(n3515), .Q(n1423) );
  XNR22 U4155 ( .A(n1472), .B(n3538), .Q(n3515) );
  NOR42 U4156 ( .A(n2800), .B(n2801), .C(n2802), .D(n2803), .Q(n2799) );
  AOI220 U4157 ( .A(n1779), .B(n6313), .C(n1142), .D(inst_out[11]), .Q(n1778)
         );
  AOI220 U4158 ( .A(n1783), .B(n6314), .C(n1142), .D(inst_out[2]), .Q(n1782)
         );
  AOI220 U4159 ( .A(n1795), .B(n6312), .C(n1142), .D(inst_out[7]), .Q(n1794)
         );
  OAI310 U4160 ( .A(n6357), .B(n6347), .C(n3564), .D(n3504), .Q(n3549) );
  NAND30 U4161 ( .A(n6513), .B(n1379), .C(n4041), .Q(n4037) );
  OAI220 U4162 ( .A(n6347), .B(n6514), .C(n1420), .D(n6517), .Q(n3556) );
  AOI220 U4163 ( .A(n6355), .B(n6193), .C(n1294), .D(n6347), .Q(n3599) );
  CLKIN6 U4164 ( .A(n1993), .Q(n6280) );
  NAND43 U4165 ( .A(n1891), .B(n1892), .C(n1893), .D(n1894), .Q(n1869) );
  NOR40 U4166 ( .A(n4333), .B(n4334), .C(n6341), .D(n4335), .Q(n4332) );
  NOR41 U4167 ( .A(n6321), .B(n4280), .C(n4281), .D(n4282), .Q(n4279) );
  AOI2112 U4168 ( .A(n6222), .B(n1381), .C(n4311), .D(n4312), .Q(n4310) );
  NOR41 U4169 ( .A(n4320), .B(n4321), .C(n4322), .D(n4323), .Q(n4319) );
  AOI222 U4170 ( .A(n4283), .B(n3625), .C(n3622), .D(n1991), .Q(n4280) );
  NOR42 U4171 ( .A(n1903), .B(n1904), .C(n1905), .D(n1906), .Q(n1892) );
  NOR22 U4172 ( .A(n6486), .B(inst_out[0]), .Q(n1839) );
  NOR42 U4173 ( .A(n3031), .B(n3032), .C(n3033), .D(n3034), .Q(n3030) );
  NOR31 U4174 ( .A(n6097), .B(n3288), .C(n3287), .Q(n3281) );
  OAI220 U4175 ( .A(n5053), .B(n6565), .C(n5052), .D(n6564), .Q(n3288) );
  NOR31 U4176 ( .A(n2149), .B(n2148), .C(n2147), .Q(n6098) );
  INV3 U4177 ( .A(n6098), .Q(n6099) );
  NAND31 U4178 ( .A(n2376), .B(n2374), .C(n2375), .Q(n6100) );
  INV3 U4179 ( .A(n6100), .Q(n6101) );
  NOR41 U4180 ( .A(n2378), .B(n2379), .C(n2380), .D(n2381), .Q(n2377) );
  NOR24 U4181 ( .A(n2912), .B(n2911), .Q(n6102) );
  NOR31 U4182 ( .A(n6103), .B(n2910), .C(n2909), .Q(n2903) );
  CLKIN6 U4183 ( .A(n6102), .Q(n6103) );
  OAI222 U4184 ( .A(n5039), .B(n6560), .C(n5038), .D(n1932), .Q(n2909) );
  OAI222 U4185 ( .A(n5035), .B(n6578), .C(n5034), .D(n1928), .Q(n2911) );
  NAND31 U4186 ( .A(n2771), .B(n2769), .C(n2770), .Q(n6104) );
  NAND23 U4187 ( .A(n2772), .B(n6105), .Q(\instruction_decode/old_data_1 [6])
         );
  INV3 U4188 ( .A(n6104), .Q(n6105) );
  NOR41 U4189 ( .A(n2773), .B(n2774), .C(n2775), .D(n2776), .Q(n2772) );
  NAND31 U4190 ( .A(n4561), .B(n4560), .C(n4562), .Q(n6106) );
  INV3 U4191 ( .A(n6106), .Q(n6107) );
  XNR21 U4192 ( .A(write_register[4]), .B(n6221), .Q(n4562) );
  NOR31 U4193 ( .A(n6109), .B(n2385), .C(n2384), .Q(n2383) );
  OAI222 U4194 ( .A(n5093), .B(n6541), .C(n5092), .D(n6536), .Q(n2386) );
  OAI222 U4195 ( .A(n5329), .B(n6550), .C(n5328), .D(n2009), .Q(n2387) );
  NOR22 U4196 ( .A(n2391), .B(n2390), .Q(n6110) );
  NOR31 U4197 ( .A(n6111), .B(n2389), .C(n2388), .Q(n2382) );
  INV3 U4198 ( .A(n6110), .Q(n6111) );
  OAI220 U4199 ( .A(n5337), .B(n6523), .C(n5336), .D(n6519), .Q(n2388) );
  OAI220 U4200 ( .A(n4975), .B(n6532), .C(n4974), .D(n6527), .Q(n2389) );
  NOR31 U4201 ( .A(n1917), .B(n1915), .C(n1916), .Q(n6112) );
  INV3 U4202 ( .A(n6112), .Q(n6113) );
  NOR31 U4203 ( .A(n2506), .B(n2504), .C(n2505), .Q(n6114) );
  INV3 U4204 ( .A(n6114), .Q(n6115) );
  NOR31 U4205 ( .A(n6117), .B(n2158), .C(n2157), .Q(n2151) );
  NOR31 U4206 ( .A(n6119), .B(n2305), .C(n2304), .Q(n2298) );
  OAI221 U4207 ( .A(n4967), .B(n6533), .C(n4966), .D(n2013), .Q(n2305) );
  NOR31 U4208 ( .A(n2569), .B(n2567), .C(n2568), .Q(n6120) );
  INV3 U4209 ( .A(n6120), .Q(n6121) );
  NAND31 U4210 ( .A(n2981), .B(n2979), .C(n2980), .Q(n6122) );
  NAND22 U4211 ( .A(n2982), .B(n6123), .Q(\instruction_decode/old_data_1 [26])
         );
  INV3 U4212 ( .A(n6122), .Q(n6123) );
  NOR41 U4213 ( .A(n2983), .B(n2984), .C(n2985), .D(n2986), .Q(n2982) );
  NOR31 U4214 ( .A(n2065), .B(n2063), .C(n2064), .Q(n6124) );
  INV3 U4215 ( .A(n6124), .Q(n6125) );
  NOR31 U4216 ( .A(n3152), .B(n3153), .C(n3151), .Q(n6126) );
  INV3 U4217 ( .A(n6126), .Q(n6127) );
  NOR33 U4218 ( .A(n6129), .B(n2242), .C(n2241), .Q(n2235) );
  CLKIN6 U4219 ( .A(n6128), .Q(n6129) );
  OAI221 U4220 ( .A(n4963), .B(n6524), .C(n4962), .D(n2015), .Q(n2241) );
  NOR31 U4221 ( .A(n6131), .B(n1935), .C(n1933), .Q(n1919) );
  NOR31 U4222 ( .A(n2589), .B(n2590), .C(n2588), .Q(n6132) );
  INV3 U4223 ( .A(n6132), .Q(n6133) );
  NOR31 U4224 ( .A(n6135), .B(n2515), .C(n2514), .Q(n2508) );
  OAI221 U4225 ( .A(n5013), .B(n6530), .C(n5012), .D(n6528), .Q(n2515) );
  NOR31 U4226 ( .A(n3174), .B(n3173), .C(n3172), .Q(n6136) );
  INV3 U4227 ( .A(n6136), .Q(n6137) );
  NOR31 U4228 ( .A(n3215), .B(n3216), .C(n3214), .Q(n6138) );
  INV3 U4229 ( .A(n6138), .Q(n6139) );
  NOR31 U4230 ( .A(n2674), .B(n2673), .C(n2672), .Q(n6140) );
  INV3 U4231 ( .A(n6140), .Q(n6141) );
  NAND31 U4232 ( .A(n3002), .B(n3000), .C(n3001), .Q(n6142) );
  INV3 U4233 ( .A(n6142), .Q(n6143) );
  NOR41 U4234 ( .A(n3004), .B(n3005), .C(n3006), .D(n3007), .Q(n3003) );
  NAND34 U4235 ( .A(n1728), .B(n4568), .C(n6145), .Q(n4423) );
  INV6 U4236 ( .A(n6144), .Q(n6145) );
  XNR22 U4237 ( .A(write_register_ex[2]), .B(rt[2]), .Q(n4567) );
  NOR32 U4238 ( .A(n4569), .B(n4570), .C(n4571), .Q(n4568) );
  NAND30 U4239 ( .A(n5734), .B(n5699), .C(n5694), .Q(n6146) );
  NAND22 U4240 ( .A(n4544), .B(n6147), .Q(n4479) );
  CLKIN2 U4241 ( .A(n6146), .Q(n6147) );
  INV2 U4242 ( .A(n4479), .Q(n1467) );
  NAND31 U4243 ( .A(n2939), .B(n2937), .C(n2938), .Q(n6148) );
  NAND24 U4244 ( .A(n2940), .B(n6149), .Q(\instruction_decode/old_data_1 [28])
         );
  INV3 U4245 ( .A(n6148), .Q(n6149) );
  NOR31 U4246 ( .A(n6151), .B(n2599), .C(n2598), .Q(n2592) );
  OAI221 U4247 ( .A(n5003), .B(n6529), .C(n5002), .D(n6527), .Q(n2599) );
  NOR31 U4248 ( .A(n6153), .B(n3183), .C(n3182), .Q(n3176) );
  OAI221 U4249 ( .A(n4981), .B(n6557), .C(n4980), .D(n6554), .Q(n3182) );
  OAI221 U4250 ( .A(n4979), .B(n6566), .C(n4978), .D(n6563), .Q(n3183) );
  NOR31 U4251 ( .A(n6155), .B(n3225), .C(n3224), .Q(n3218) );
  OAI220 U4252 ( .A(n5071), .B(n6566), .C(n5070), .D(n1930), .Q(n3225) );
  NOR31 U4253 ( .A(n2733), .B(n2732), .C(n2731), .Q(n6156) );
  INV3 U4254 ( .A(n6156), .Q(n6157) );
  NOR31 U4255 ( .A(n2000), .B(n1999), .C(n1998), .Q(n6158) );
  INV3 U4256 ( .A(n6158), .Q(n6159) );
  NOR31 U4257 ( .A(n6161), .B(n2683), .C(n2682), .Q(n2676) );
  OAI221 U4258 ( .A(n4951), .B(n6529), .C(n4950), .D(n6527), .Q(n2683) );
  NAND31 U4259 ( .A(n2855), .B(n2853), .C(n2854), .Q(n6162) );
  INV3 U4260 ( .A(n6162), .Q(n6163) );
  NOR31 U4261 ( .A(n3257), .B(n3258), .C(n3256), .Q(n6164) );
  INV3 U4262 ( .A(n6164), .Q(n6165) );
  NOR31 U4263 ( .A(n2128), .B(n2127), .C(n2126), .Q(n6166) );
  INV3 U4264 ( .A(n6166), .Q(n6167) );
  NOR31 U4265 ( .A(n2211), .B(n2212), .C(n2210), .Q(n6168) );
  NOR23 U4266 ( .A(n6169), .B(n2213), .Q(n2209) );
  INV3 U4267 ( .A(n6168), .Q(n6169) );
  NAND22 U4268 ( .A(n3672), .B(n3668), .Q(n6170) );
  NAND24 U4269 ( .A(n3673), .B(n6171), .Q(n3633) );
  INV3 U4270 ( .A(n6170), .Q(n6171) );
  NOR22 U4271 ( .A(n3744), .B(n1407), .Q(n3673) );
  NOR31 U4272 ( .A(n3631), .B(n3633), .C(n3632), .Q(n6218) );
  INV3 U4273 ( .A(n3633), .Q(n6214) );
  NOR31 U4274 ( .A(n6173), .B(n2741), .C(n2742), .Q(n2735) );
  OAI221 U4275 ( .A(n5127), .B(n6562), .C(n5126), .D(n1932), .Q(n2741) );
  NOR31 U4276 ( .A(n6175), .B(n2017), .C(n2016), .Q(n2002) );
  OAI221 U4277 ( .A(n5049), .B(n6535), .C(n5048), .D(n6527), .Q(n2017) );
  CLKIN1 U4278 ( .A(n1472), .Q(n6176) );
  NOR23 U4279 ( .A(n4170), .B(n4171), .Q(n4062) );
  NOR31 U4280 ( .A(n6180), .B(n3267), .C(n3266), .Q(n3260) );
  OAI221 U4281 ( .A(n5313), .B(n6556), .C(n5312), .D(n6554), .Q(n3266) );
  OAI221 U4282 ( .A(n4971), .B(n6565), .C(n4970), .D(n1930), .Q(n3267) );
  NOR31 U4283 ( .A(n2464), .B(n2462), .C(n2463), .Q(n6181) );
  INV3 U4284 ( .A(n6181), .Q(n6182) );
  NOR31 U4285 ( .A(n3110), .B(n3111), .C(n3109), .Q(n6183) );
  INV3 U4286 ( .A(n6183), .Q(n6184) );
  NOR31 U4287 ( .A(n6186), .B(n2137), .C(n2136), .Q(n2130) );
  OAI221 U4288 ( .A(n5159), .B(n6534), .C(n5158), .D(n6528), .Q(n2137) );
  NOR31 U4289 ( .A(n3047), .B(n3048), .C(n3046), .Q(n6187) );
  INV3 U4290 ( .A(n6187), .Q(n6188) );
  NOR31 U4291 ( .A(n2922), .B(n2920), .C(n2921), .Q(n6189) );
  NOR24 U4292 ( .A(n6190), .B(n2923), .Q(n2919) );
  INV3 U4293 ( .A(n6189), .Q(n6190) );
  NOR31 U4294 ( .A(n2838), .B(n2837), .C(n2836), .Q(n6191) );
  INV3 U4295 ( .A(n6191), .Q(n6192) );
  NAND31 U4296 ( .A(n2897), .B(n2895), .C(n2896), .Q(n6196) );
  NAND22 U4297 ( .A(n2898), .B(n6197), .Q(\instruction_decode/old_data_1 [2])
         );
  INV3 U4298 ( .A(n6196), .Q(n6197) );
  NOR41 U4299 ( .A(n2899), .B(n2900), .C(n2901), .D(n2902), .Q(n2898) );
  OAI222 U4300 ( .A(n4961), .B(n6569), .C(n4960), .D(n6563), .Q(n2931) );
  NOR42 U4301 ( .A(n2441), .B(n2442), .C(n2443), .D(n2444), .Q(n2440) );
  OAI222 U4302 ( .A(n5195), .B(n6578), .C(n5194), .D(n6572), .Q(n2907) );
  NOR41 U4303 ( .A(n2300), .B(n2301), .C(n2302), .D(n2303), .Q(n2299) );
  NOR41 U4304 ( .A(n2451), .B(n2452), .C(n2453), .D(n2454), .Q(n2445) );
  OAI222 U4305 ( .A(n5243), .B(n6570), .C(n5242), .D(n6563), .Q(n2864) );
  NAND43 U4306 ( .A(n2164), .B(n2165), .C(n2166), .D(n2167), .Q(
        \instruction_decode/old_data_2 [31]) );
  NOR42 U4307 ( .A(n2105), .B(n2106), .C(n2107), .D(n2108), .Q(n2104) );
  OAI222 U4308 ( .A(n4963), .B(n6560), .C(n4962), .D(n1932), .Q(n2930) );
  NOR41 U4309 ( .A(n2283), .B(n2284), .C(n2285), .D(n2286), .Q(n2277) );
  NAND43 U4310 ( .A(n2248), .B(n2249), .C(n2250), .D(n2251), .Q(
        \instruction_decode/old_data_2 [28]) );
  NAND43 U4311 ( .A(n3084), .B(n3085), .C(n3086), .D(n3087), .Q(
        \instruction_decode/old_data_1 [21]) );
  NOR42 U4312 ( .A(n3088), .B(n3089), .C(n3090), .D(n3091), .Q(n3087) );
  NOR41 U4313 ( .A(n2115), .B(n2116), .C(n2117), .D(n2118), .Q(n2109) );
  NAND43 U4314 ( .A(n3336), .B(n3337), .C(n3338), .D(n3339), .Q(
        \instruction_decode/old_data_1 [0]) );
  NOR41 U4315 ( .A(n2346), .B(n2347), .C(n2348), .D(n2349), .Q(n2340) );
  NOR41 U4316 ( .A(n2720), .B(n2721), .C(n2722), .D(n2723), .Q(n2714) );
  NAND43 U4317 ( .A(n2080), .B(n2081), .C(n2082), .D(n2083), .Q(
        \instruction_decode/old_data_2 [6]) );
  NOR42 U4318 ( .A(n2084), .B(n2085), .C(n2086), .D(n2087), .Q(n2083) );
  NAND43 U4319 ( .A(n2416), .B(n2417), .C(n2418), .D(n2419), .Q(
        \instruction_decode/old_data_2 [20]) );
  NOR41 U4320 ( .A(n3098), .B(n3099), .C(n3100), .D(n3101), .Q(n3092) );
  XOR22 U4321 ( .A(\instruction_decode/old_data_1 [30]), .B(
        \instruction_decode/old_data_2 [30]), .Q(n1907) );
  AOI221 U4322 ( .A(n6332), .B(data_2[2]), .C(n5815), .D(ram_adr[2]), .Q(n4435) );
  NOR42 U4323 ( .A(n2195), .B(n2196), .C(n2197), .D(n2198), .Q(n2194) );
  NOR41 U4324 ( .A(n3350), .B(n3351), .C(n3352), .D(n3353), .Q(n3344) );
  NOR41 U4325 ( .A(n3329), .B(n3330), .C(n3331), .D(n3332), .Q(n3323) );
  NAND43 U4326 ( .A(n2811), .B(n2812), .C(n2813), .D(n2814), .Q(
        \instruction_decode/old_data_1 [4]) );
  NOR42 U4327 ( .A(n2815), .B(n2816), .C(n2817), .D(n2818), .Q(n2814) );
  NAND43 U4328 ( .A(n3063), .B(n3064), .C(n3065), .D(n3066), .Q(
        \instruction_decode/old_data_1 [22]) );
  NOR42 U4329 ( .A(n3067), .B(n3068), .C(n3069), .D(n3070), .Q(n3066) );
  NOR41 U4330 ( .A(n2094), .B(n2095), .C(n2096), .D(n2097), .Q(n2088) );
  INV2 U4331 ( .A(n6202), .Q(n6203) );
  NOR41 U4332 ( .A(n2825), .B(n2826), .C(n2827), .D(n2828), .Q(n2819) );
  NAND43 U4333 ( .A(n2647), .B(n2648), .C(n2649), .D(n2650), .Q(
        \instruction_decode/old_data_2 [10]) );
  NOR41 U4334 ( .A(n3077), .B(n3078), .C(n3079), .D(n3080), .Q(n3071) );
  NOR42 U4335 ( .A(n2315), .B(n2316), .C(n2317), .D(n2318), .Q(n2314) );
  NAND22 U4336 ( .A(n4238), .B(n3436), .Q(n3443) );
  NAND43 U4337 ( .A(n2227), .B(n2228), .C(n2229), .D(n2230), .Q(
        \instruction_decode/old_data_2 [29]) );
  NAND22 U4338 ( .A(n6321), .B(n1420), .Q(n6243) );
  OAI221 U4339 ( .A(n4895), .B(n6588), .C(n4894), .D(n1926), .Q(n2950) );
  OAI221 U4340 ( .A(n4935), .B(n6589), .C(n4934), .D(n1926), .Q(n2866) );
  CLKIN6 U4341 ( .A(n4404), .Q(n6505) );
  NOR41 U4342 ( .A(n2325), .B(n2326), .C(n2327), .D(n2328), .Q(n2319) );
  OAI221 U4343 ( .A(n4983), .B(n6578), .C(n4982), .D(n6573), .Q(n2953) );
  OAI221 U4344 ( .A(n5099), .B(n6579), .C(n5098), .D(n1928), .Q(n2869) );
  NAND43 U4345 ( .A(n2395), .B(n2396), .C(n2397), .D(n2398), .Q(
        \instruction_decode/old_data_2 [21]) );
  OAI222 U4346 ( .A(n1425), .B(n1360), .C(n4326), .D(n4327), .Q(n4324) );
  NAND43 U4347 ( .A(n2958), .B(n2959), .C(n2960), .D(n2961), .Q(
        \instruction_decode/old_data_1 [27]) );
  NAND43 U4348 ( .A(n2790), .B(n2791), .C(n2792), .D(n2793), .Q(
        \instruction_decode/old_data_1 [5]) );
  NOR42 U4349 ( .A(n2794), .B(n2795), .C(n2796), .D(n2797), .Q(n2793) );
  NOR41 U4350 ( .A(n3140), .B(n3141), .C(n3142), .D(n3143), .Q(n3134) );
  NAND43 U4351 ( .A(n3021), .B(n3022), .C(n3023), .D(n3024), .Q(
        \instruction_decode/old_data_1 [24]) );
  NOR42 U4352 ( .A(n3025), .B(n3026), .C(n3027), .D(n3028), .Q(n3024) );
  XNR22 U4353 ( .A(write_register_ex[0]), .B(rt[0]), .Q(n4566) );
  NOR41 U4354 ( .A(n2972), .B(n2973), .C(n2974), .D(n2975), .Q(n2966) );
  NOR41 U4355 ( .A(n2804), .B(n2805), .C(n2806), .D(n2807), .Q(n2798) );
  NOR41 U4356 ( .A(n3035), .B(n3036), .C(n3037), .D(n3038), .Q(n3029) );
  NOR21 U4357 ( .A(n4130), .B(n1372), .Q(n4061) );
  INV3 U4358 ( .A(n3966), .Q(n1387) );
  OAI222 U4359 ( .A(n4853), .B(n6589), .C(n4852), .D(n1926), .Q(n2887) );
  OAI221 U4360 ( .A(n4871), .B(n6588), .C(n4870), .D(n1926), .Q(n2929) );
  OAI221 U4361 ( .A(n4959), .B(n6578), .C(n4958), .D(n1928), .Q(n2932) );
  NOR41 U4362 ( .A(n3014), .B(n3015), .C(n3016), .D(n3017), .Q(n3008) );
  OAI221 U4363 ( .A(n4985), .B(n6569), .C(n4984), .D(n1930), .Q(n2952) );
  OAI221 U4364 ( .A(n5351), .B(n6560), .C(n5350), .D(n6555), .Q(n2951) );
  OAI221 U4365 ( .A(n5241), .B(n6579), .C(n5240), .D(n6573), .Q(n2865) );
  OAI221 U4366 ( .A(n5101), .B(n6570), .C(n5100), .D(n6563), .Q(n2868) );
  OAI221 U4367 ( .A(n5103), .B(n6561), .C(n5102), .D(n1932), .Q(n2867) );
  NOR42 U4368 ( .A(n2174), .B(n2175), .C(n2176), .D(n2177), .Q(n2173) );
  CLKIN3 U4369 ( .A(n3973), .Q(n1446) );
  NOR42 U4370 ( .A(n2941), .B(n2942), .C(n2943), .D(n2944), .Q(n2940) );
  OAI221 U4371 ( .A(n5037), .B(n6569), .C(n5036), .D(n6563), .Q(n2910) );
  NOR20 U4372 ( .A(n3527), .B(n3528), .Q(n3516) );
  NOR22 U4373 ( .A(n3564), .B(n3562), .Q(n3528) );
  NOR41 U4374 ( .A(n1883), .B(n1884), .C(n1885), .D(n1886), .Q(n1872) );
  NOR42 U4375 ( .A(n1887), .B(n1888), .C(n1889), .D(n1890), .Q(n1871) );
  NOR42 U4376 ( .A(n1907), .B(n1908), .C(n1909), .D(n1910), .Q(n1891) );
  NOR41 U4377 ( .A(n2867), .B(n2868), .C(n2869), .D(n2870), .Q(n2861) );
  NOR42 U4378 ( .A(n2258), .B(n2259), .C(n2260), .D(n2261), .Q(n2257) );
  OAI221 U4379 ( .A(n5117), .B(n6578), .C(n5116), .D(n6572), .Q(n2949) );
  NOR41 U4380 ( .A(n2783), .B(n2784), .C(n2785), .D(n2786), .Q(n2777) );
  NOR41 U4381 ( .A(n2951), .B(n2952), .C(n2953), .D(n2954), .Q(n2945) );
  XOR22 U4382 ( .A(\instruction_decode/old_data_1 [11]), .B(
        \instruction_decode/old_data_2 [11]), .Q(n1878) );
  NAND42 U4383 ( .A(n3294), .B(n3295), .C(n3296), .D(n3297), .Q(
        \instruction_decode/old_data_1 [11]) );
  INV2 U4384 ( .A(n4335), .Q(n1318) );
  OAI221 U4385 ( .A(n1416), .B(n1320), .C(n6349), .D(n1338), .Q(n4335) );
  NOR42 U4386 ( .A(n2884), .B(n2885), .C(n2886), .D(n2887), .Q(n2883) );
  NAND42 U4387 ( .A(n2626), .B(n2627), .C(n2628), .D(n2629), .Q(
        \instruction_decode/old_data_2 [11]) );
  OAI2111 U4388 ( .A(n1420), .B(n3564), .C(n4330), .D(n4331), .Q(n4329) );
  AOI310 U4389 ( .A(n1310), .B(n1415), .C(n1318), .D(n4332), .Q(n4331) );
  XOR22 U4390 ( .A(\instruction_decode/old_data_1 [12]), .B(
        \instruction_decode/old_data_2 [12]), .Q(n1877) );
  NAND42 U4391 ( .A(n3273), .B(n3274), .C(n3275), .D(n3276), .Q(
        \instruction_decode/old_data_1 [12]) );
  INV3 U4392 ( .A(n3811), .Q(n1401) );
  NAND42 U4393 ( .A(n2605), .B(n2606), .C(n2607), .D(n2608), .Q(
        \instruction_decode/old_data_2 [12]) );
  XOR22 U4394 ( .A(\instruction_decode/old_data_1 [15]), .B(
        \instruction_decode/old_data_2 [15]), .Q(n1898) );
  NAND42 U4395 ( .A(n3231), .B(n3232), .C(n3233), .D(n3234), .Q(
        \instruction_decode/old_data_1 [15]) );
  NOR41 U4396 ( .A(n3304), .B(n3305), .C(n3306), .D(n3307), .Q(n3303) );
  XOR22 U4397 ( .A(\instruction_decode/old_data_1 [14]), .B(
        \instruction_decode/old_data_2 [14]), .Q(n1875) );
  NAND42 U4398 ( .A(n1911), .B(n1912), .C(n1913), .D(n1914), .Q(
        \instruction_decode/reg_MAPP/n3641 ) );
  NAND42 U4399 ( .A(n2563), .B(n2564), .C(n2565), .D(n2566), .Q(
        \instruction_decode/old_data_2 [14]) );
  XOR22 U4400 ( .A(\instruction_decode/old_data_1 [7]), .B(
        \instruction_decode/old_data_2 [7]), .Q(n1882) );
  NAND42 U4401 ( .A(n2748), .B(n2749), .C(n2750), .D(n2751), .Q(
        \instruction_decode/old_data_1 [7]) );
  NOR41 U4402 ( .A(n2636), .B(n2637), .C(n2638), .D(n2639), .Q(n2635) );
  XOR22 U4403 ( .A(\instruction_decode/old_data_1 [23]), .B(
        \instruction_decode/old_data_2 [23]), .Q(n1906) );
  INV3 U4404 ( .A(n3718), .Q(n1410) );
  NOR22 U4405 ( .A(n5945), .B(n1772), .Q(n1985) );
  NAND26 U4406 ( .A(n1768), .B(n6249), .Q(n1772) );
  OAI210 U4407 ( .A(n1408), .B(n3737), .C(n3740), .Q(n3762) );
  CLKIN6 U4408 ( .A(n3439), .Q(n6198) );
  NOR41 U4409 ( .A(n3283), .B(n3284), .C(n3285), .D(n3286), .Q(n3282) );
  NAND42 U4410 ( .A(n2143), .B(n2144), .C(n2145), .D(n2146), .Q(
        \instruction_decode/old_data_2 [3]) );
  NAND22 U4411 ( .A(n3910), .B(n1393), .Q(n3899) );
  INV3 U4412 ( .A(n3907), .Q(n1393) );
  XOR22 U4413 ( .A(\instruction_decode/old_data_1 [19]), .B(
        \instruction_decode/old_data_2 [19]), .Q(n1902) );
  NOR41 U4414 ( .A(n2615), .B(n2616), .C(n2617), .D(n2618), .Q(n2614) );
  CLKBU12 U4415 ( .A(n3691), .Q(n6204) );
  NAND42 U4416 ( .A(n2542), .B(n2543), .C(n2544), .D(n2545), .Q(
        \instruction_decode/old_data_2 [15]) );
  XOR22 U4417 ( .A(\instruction_decode/old_data_1 [16]), .B(
        \instruction_decode/old_data_2 [16]), .Q(n1897) );
  AOI211 U4418 ( .A(n3564), .B(n1420), .C(n4328), .Q(n4326) );
  NOR41 U4419 ( .A(n3241), .B(n3242), .C(n3243), .D(n3244), .Q(n3240) );
  XOR22 U4420 ( .A(\instruction_decode/old_data_1 [0]), .B(
        \instruction_decode/old_data_2 [0]), .Q(n1890) );
  NAND22 U4421 ( .A(n1455), .B(n3777), .Q(n3742) );
  CLKIN1 U4422 ( .A(n3786), .Q(n1455) );
  XOR22 U4423 ( .A(\instruction_decode/old_data_1 [8]), .B(
        \instruction_decode/old_data_2 [8]), .Q(n1881) );
  NAND42 U4424 ( .A(n2521), .B(n2522), .C(n2523), .D(n2524), .Q(
        \instruction_decode/old_data_2 [16]) );
  XOR22 U4425 ( .A(\instruction_decode/old_data_1 [2]), .B(
        \instruction_decode/old_data_2 [2]), .Q(n1887) );
  NAND42 U4426 ( .A(n2059), .B(n2060), .C(n2061), .D(n2062), .Q(
        \instruction_decode/old_data_2 [7]) );
  NAND21 U4427 ( .A(n3691), .B(n3692), .Q(n3690) );
  XOR22 U4428 ( .A(\instruction_decode/old_data_1 [3]), .B(
        \instruction_decode/old_data_2 [3]), .Q(n1886) );
  XOR22 U4429 ( .A(\instruction_decode/old_data_1 [17]), .B(
        \instruction_decode/old_data_2 [17]), .Q(n1896) );
  XOR22 U4430 ( .A(\instruction_decode/old_data_1 [20]), .B(
        \instruction_decode/old_data_2 [20]), .Q(n1901) );
  NOR41 U4431 ( .A(n2758), .B(n2759), .C(n2760), .D(n2761), .Q(n2757) );
  XOR22 U4432 ( .A(\instruction_decode/old_data_1 [24]), .B(
        \instruction_decode/old_data_2 [24]), .Q(n1905) );
  XOR22 U4433 ( .A(\instruction_decode/old_data_2 [18]), .B(
        \instruction_decode/old_data_1 [18]), .Q(n1895) );
  NAND42 U4434 ( .A(n2500), .B(n2501), .C(n2502), .D(n2503), .Q(
        \instruction_decode/old_data_2 [17]) );
  XOR22 U4435 ( .A(\instruction_decode/old_data_1 [9]), .B(
        \instruction_decode/old_data_2 [9]), .Q(n1880) );
  XOR22 U4436 ( .A(\instruction_decode/old_data_1 [27]), .B(
        \instruction_decode/old_data_2 [27]), .Q(n1910) );
  XOR22 U4437 ( .A(\instruction_decode/old_data_1 [10]), .B(
        \instruction_decode/old_data_2 [10]), .Q(n1879) );
  NAND22 U4438 ( .A(n3471), .B(n6250), .Q(n4242) );
  XNR22 U4439 ( .A(n1472), .B(n1425), .Q(n3471) );
  XOR22 U4440 ( .A(\instruction_decode/old_data_1 [1]), .B(
        \instruction_decode/old_data_2 [1]), .Q(n1889) );
  XOR22 U4441 ( .A(\instruction_decode/old_data_1 [21]), .B(
        \instruction_decode/old_data_2 [21]), .Q(n1900) );
  XOR22 U4442 ( .A(\instruction_decode/old_data_1 [25]), .B(
        \instruction_decode/old_data_2 [25]), .Q(n1904) );
  NAND43 U4443 ( .A(n2290), .B(n2291), .C(n2292), .D(n2293), .Q(
        \instruction_decode/old_data_2 [26]) );
  XOR22 U4444 ( .A(\instruction_decode/old_data_1 [4]), .B(
        \instruction_decode/old_data_2 [4]), .Q(n1885) );
  NOR41 U4445 ( .A(n2552), .B(n2553), .C(n2554), .D(n2555), .Q(n2551) );
  XOR22 U4446 ( .A(\instruction_decode/old_data_1 [22]), .B(
        \instruction_decode/old_data_2 [22]), .Q(n1899) );
  NOR41 U4447 ( .A(n2363), .B(n2364), .C(n2365), .D(n2366), .Q(n2362) );
  NOR41 U4448 ( .A(n2342), .B(n2343), .C(n2344), .D(n2345), .Q(n2341) );
  NOR41 U4449 ( .A(n2531), .B(n2532), .C(n2533), .D(n2534), .Q(n2530) );
  XOR22 U4450 ( .A(\instruction_decode/old_data_1 [5]), .B(
        \instruction_decode/old_data_2 [5]), .Q(n1884) );
  OAI2112 U4451 ( .A(n5699), .B(n5733), .C(n4405), .D(n1481), .Q(n3627) );
  NOR41 U4452 ( .A(n3199), .B(n3200), .C(n3201), .D(n3202), .Q(n3198) );
  XOR22 U4453 ( .A(\instruction_decode/old_data_1 [6]), .B(
        \instruction_decode/old_data_2 [6]), .Q(n1883) );
  NOR41 U4454 ( .A(n2489), .B(n2490), .C(n2491), .D(n2492), .Q(n2488) );
  NOR41 U4455 ( .A(n2716), .B(n2717), .C(n2718), .D(n2719), .Q(n2715) );
  NOR41 U4456 ( .A(n2048), .B(n2049), .C(n2050), .D(n2051), .Q(n2047) );
  NOR41 U4457 ( .A(n2821), .B(n2822), .C(n2823), .D(n2824), .Q(n2820) );
  NOR41 U4458 ( .A(n2426), .B(n2427), .C(n2428), .D(n2429), .Q(n2425) );
  NOR22 U4459 ( .A(n6238), .B(n1468), .Q(n4427) );
  NOR41 U4460 ( .A(n2111), .B(n2112), .C(n2113), .D(n2114), .Q(n2110) );
  NOR21 U4461 ( .A(n3436), .B(n4238), .Q(n3442) );
  XNR22 U4462 ( .A(n1472), .B(n6199), .Q(n4238) );
  NOR41 U4463 ( .A(n2090), .B(n2091), .C(n2092), .D(n2093), .Q(n2089) );
  XNR22 U4464 ( .A(n1472), .B(n4227), .Q(n4175) );
  INV2 U4465 ( .A(n6237), .Q(n6238) );
  NOR41 U4466 ( .A(n2405), .B(n2406), .C(n2407), .D(n2408), .Q(n2404) );
  NOR41 U4467 ( .A(n2657), .B(n2658), .C(n2659), .D(n2660), .Q(n2656) );
  NOR41 U4468 ( .A(n2779), .B(n2780), .C(n2781), .D(n2782), .Q(n2778) );
  OAI2112 U4469 ( .A(n4050), .B(n4051), .C(n4052), .D(n4044), .Q(n4049) );
  NAND22 U4470 ( .A(n1377), .B(n6261), .Q(n4044) );
  XNR21 U4471 ( .A(n3870), .B(n6322), .Q(n3851) );
  OAI212 U4472 ( .A(n1356), .B(n1423), .C(n3563), .Q(n4241) );
  AOI2112 U4473 ( .A(n4058), .B(n4059), .C(n4060), .D(n4061), .Q(n4056) );
  AOI221 U4474 ( .A(n6332), .B(data_2[14]), .C(n5815), .D(ram_adr[14]), .Q(
        n4453) );
  NAND22 U4475 ( .A(n4110), .B(n4111), .Q(n4057) );
  XNR21 U4476 ( .A(n6321), .B(n1436), .Q(n4110) );
  NOR20 U4477 ( .A(n1369), .B(n1371), .Q(n6200) );
  INV3 U4478 ( .A(n6200), .Q(n6201) );
  NOR21 U4479 ( .A(n1486), .B(n1468), .Q(n6202) );
  NOR20 U4480 ( .A(n6203), .B(n1484), .Q(n6327) );
  INV10 U4481 ( .A(n4423), .Q(n1486) );
  NAND22 U4482 ( .A(n3832), .B(n6205), .Q(n6206) );
  NAND24 U4483 ( .A(n6206), .B(n1392), .Q(n3639) );
  INV0 U4484 ( .A(n3827), .Q(n6205) );
  INV3 U4485 ( .A(n3832), .Q(n1398) );
  NAND22 U4486 ( .A(n1449), .B(n6321), .Q(n6207) );
  NOR22 U4487 ( .A(n1395), .B(n3875), .Q(n3873) );
  BUF2 U4488 ( .A(n6067), .Q(n6209) );
  NAND22 U4489 ( .A(n6321), .B(n6345), .Q(n6211) );
  NAND26 U4490 ( .A(n6350), .B(n6210), .Q(n6212) );
  NAND28 U4491 ( .A(n6211), .B(n6212), .Q(n4165) );
  NAND31 U4492 ( .A(n3971), .B(n6213), .C(n6214), .Q(n6215) );
  NAND22 U4493 ( .A(n6215), .B(n3643), .Q(n3628) );
  NAND33 U4494 ( .A(n3641), .B(n3640), .C(n3805), .Q(n3632) );
  NAND22 U4495 ( .A(n3786), .B(n1405), .Q(n3741) );
  NOR24 U4496 ( .A(n6219), .B(n3634), .Q(n3630) );
  OAI211 U4497 ( .A(n4048), .B(n4080), .C(n4057), .Q(n4077) );
  INV1 U4498 ( .A(n4048), .Q(n1375) );
  NAND21 U4499 ( .A(n4039), .B(n6350), .Q(n6223) );
  NAND26 U4500 ( .A(n6223), .B(n6224), .Q(n3976) );
  AOI2111 U4501 ( .A(n1381), .B(n3976), .C(n1382), .D(n3974), .Q(n3913) );
  OAI210 U4502 ( .A(n3976), .B(n4037), .C(n4040), .Q(n4035) );
  NAND21 U4503 ( .A(n1472), .B(n1416), .Q(n6229) );
  NAND24 U4504 ( .A(n6350), .B(n6228), .Q(n6230) );
  NAND24 U4505 ( .A(n6229), .B(n6230), .Q(n4248) );
  CLKIN6 U4506 ( .A(n1416), .Q(n6228) );
  BUF4 U4507 ( .A(n1472), .Q(n6321) );
  NOR22 U4508 ( .A(n4248), .B(n1320), .Q(n3591) );
  NAND22 U4509 ( .A(n6234), .B(n6256), .Q(n6235) );
  INV3 U4510 ( .A(n4350), .Q(n6234) );
  CLKIN3 U4511 ( .A(\execute/op_21 [14]), .Q(n1437) );
  OAI221 U4512 ( .A(n5097), .B(n6523), .C(n5096), .D(n6519), .Q(n2384) );
  NAND24 U4513 ( .A(n5734), .B(n6252), .Q(n4288) );
  NAND34 U4514 ( .A(n4413), .B(n5999), .C(n5700), .Q(n6251) );
  OAI221 U4515 ( .A(n5161), .B(n6541), .C(n5160), .D(n6537), .Q(n2407) );
  OAI221 U4516 ( .A(n5217), .B(n6540), .C(n5216), .D(n6536), .Q(n2428) );
  OAI221 U4517 ( .A(n4911), .B(n6550), .C(n4910), .D(n6545), .Q(n2408) );
  OAI221 U4518 ( .A(n4927), .B(n6549), .C(n4926), .D(n6546), .Q(n2429) );
  OAI221 U4519 ( .A(n5265), .B(n6539), .C(n5264), .D(n6536), .Q(n2554) );
  OAI221 U4520 ( .A(n5007), .B(n6540), .C(n5006), .D(n6536), .Q(n2411) );
  OAI221 U4521 ( .A(n4973), .B(n6541), .C(n4972), .D(n6537), .Q(n2390) );
  OAI221 U4522 ( .A(n5063), .B(n6540), .C(n5062), .D(n6536), .Q(n2432) );
  OAI221 U4523 ( .A(n4943), .B(n6548), .C(n4942), .D(n6545), .Q(n2555) );
  OAI221 U4524 ( .A(n5259), .B(n6540), .C(n5258), .D(n6536), .Q(n2470) );
  OAI221 U4525 ( .A(n5139), .B(n6539), .C(n5138), .D(n2011), .Q(n2558) );
  OAI221 U4526 ( .A(n4941), .B(n6549), .C(n4940), .D(n2009), .Q(n2471) );
  OAI221 U4527 ( .A(n5229), .B(n6541), .C(n5228), .D(n2011), .Q(n2365) );
  OAI221 U4528 ( .A(n5133), .B(n6540), .C(n5132), .D(n6536), .Q(n2474) );
  OAI221 U4529 ( .A(n4931), .B(n6550), .C(n4930), .D(n2009), .Q(n2366) );
  OAI221 U4530 ( .A(n5075), .B(n6541), .C(n5074), .D(n6536), .Q(n2369) );
  OAI221 U4531 ( .A(n5095), .B(n6532), .C(n5094), .D(n6527), .Q(n2385) );
  OAI221 U4532 ( .A(n5219), .B(n6531), .C(n5218), .D(n6528), .Q(n2427) );
  OAI221 U4533 ( .A(n5267), .B(n6530), .C(n5266), .D(n6528), .Q(n2553) );
  OAI221 U4534 ( .A(n5065), .B(n6531), .C(n5064), .D(n6528), .Q(n2431) );
  OAI221 U4535 ( .A(n5261), .B(n6531), .C(n5260), .D(n6528), .Q(n2469) );
  OAI221 U4536 ( .A(n5141), .B(n6530), .C(n5140), .D(n6527), .Q(n2557) );
  OAI221 U4537 ( .A(n5231), .B(n6532), .C(n5230), .D(n6528), .Q(n2364) );
  OAI221 U4538 ( .A(n5135), .B(n6531), .C(n5134), .D(n6528), .Q(n2473) );
  OAI221 U4539 ( .A(n5077), .B(n6532), .C(n5076), .D(n2013), .Q(n2368) );
  OAI221 U4540 ( .A(n5149), .B(n6520), .C(n5148), .D(n6518), .Q(n2657) );
  OAI221 U4541 ( .A(n5165), .B(n6523), .C(n5164), .D(n2015), .Q(n2405) );
  OAI221 U4542 ( .A(n5221), .B(n6522), .C(n5220), .D(n6519), .Q(n2426) );
  OAI221 U4543 ( .A(n5349), .B(n6520), .C(n5348), .D(n6518), .Q(n2661) );
  OAI221 U4544 ( .A(n5269), .B(n6521), .C(n5268), .D(n6519), .Q(n2552) );
  OAI221 U4545 ( .A(n5067), .B(n6522), .C(n5066), .D(n6519), .Q(n2430) );
  OAI221 U4546 ( .A(n5263), .B(n6522), .C(n5262), .D(n6519), .Q(n2468) );
  OAI221 U4547 ( .A(n5143), .B(n6521), .C(n5142), .D(n6518), .Q(n2556) );
  OAI221 U4548 ( .A(n5233), .B(n6523), .C(n5232), .D(n6518), .Q(n2363) );
  OAI221 U4549 ( .A(n5137), .B(n6522), .C(n5136), .D(n6519), .Q(n2472) );
  OAI221 U4550 ( .A(n5079), .B(n6523), .C(n5078), .D(n6519), .Q(n2367) );
  OAI221 U4551 ( .A(n5275), .B(n6544), .C(n5274), .D(n6537), .Q(n2071) );
  OAI221 U4552 ( .A(n4947), .B(n6553), .C(n4946), .D(n6546), .Q(n2072) );
  OAI221 U4553 ( .A(n5177), .B(n6544), .C(n5176), .D(n6537), .Q(n2075) );
  OAI221 U4554 ( .A(n5277), .B(n6535), .C(n5276), .D(n6527), .Q(n2070) );
  OAI221 U4555 ( .A(n5179), .B(n6535), .C(n5178), .D(n6527), .Q(n2074) );
  OAI221 U4556 ( .A(n5257), .B(n6526), .C(n5256), .D(n2015), .Q(n2048) );
  OAI221 U4557 ( .A(n5279), .B(n6526), .C(n5278), .D(n6519), .Q(n2069) );
  OAI221 U4558 ( .A(n5127), .B(n6526), .C(n5126), .D(n2015), .Q(n2052) );
  OAI221 U4559 ( .A(n5181), .B(n6526), .C(n5180), .D(n6518), .Q(n2073) );
  OAI221 U4560 ( .A(n4595), .B(n6415), .C(n4594), .D(n6417), .Q(n2942) );
  OAI221 U4561 ( .A(n4591), .B(n1939), .C(n4590), .D(n1940), .Q(n2921) );
  AOI220 U4562 ( .A(n6408), .B(n5427), .C(n6413), .D(n5424), .Q(n3186) );
  NOR21 U4563 ( .A(n1409), .B(n3726), .Q(n3724) );
  INV3 U4564 ( .A(\execute/op_21 [16]), .Q(n6254) );
  OAI221 U4565 ( .A(n4587), .B(n6415), .C(n4586), .D(n6417), .Q(n2879) );
  NAND21 U4566 ( .A(n1338), .B(n1417), .Q(n4247) );
  NAND21 U4567 ( .A(n1484), .B(n6267), .Q(n4425) );
  CLKIN1 U4568 ( .A(n3467), .Q(n1360) );
  NAND43 U4569 ( .A(n2185), .B(n2186), .C(n2187), .D(n2188), .Q(
        \instruction_decode/old_data_2 [30]) );
  NOR20 U4570 ( .A(n1486), .B(n1484), .Q(n6237) );
  CLKIN3 U4571 ( .A(n3874), .Q(n1394) );
  NAND22 U4572 ( .A(n6350), .B(n6347), .Q(n6244) );
  NAND22 U4573 ( .A(n6243), .B(n6244), .Q(n3562) );
  AOI221 U4574 ( .A(n4297), .B(n4298), .C(n3757), .D(n3755), .Q(n4296) );
  AOI221 U4575 ( .A(n4294), .B(n4295), .C(n3718), .D(n3716), .Q(n4293) );
  INV6 U4576 ( .A(n3692), .Q(n1310) );
  NOR21 U4577 ( .A(n5942), .B(n6254), .Q(n6253) );
  INV2 U4578 ( .A(n3888), .Q(n1395) );
  AOI222 U4579 ( .A(n6330), .B(data_2[1]), .C(ram_adr[1]), .D(n5816), .Q(n4447) );
  AOI220 U4580 ( .A(n6329), .B(data_2[11]), .C(n5816), .D(ram_adr[11]), .Q(
        n4456) );
  CLKIN6 U4581 ( .A(rt[0]), .Q(n1485) );
  NAND21 U4582 ( .A(n5700), .B(n5734), .Q(n6239) );
  NAND33 U4583 ( .A(n4413), .B(n5999), .C(n6240), .Q(n6267) );
  NOR24 U4584 ( .A(n5733), .B(n5732), .Q(n4413) );
  INV2 U4585 ( .A(n5942), .Q(n6489) );
  XNR22 U4586 ( .A(n1472), .B(n4236), .Q(n3419) );
  AOI211 U4587 ( .A(n3848), .B(n3849), .C(n3846), .Q(n3847) );
  CLKIN4 U4588 ( .A(n6948), .Q(n6947) );
  CLKIN6 U4589 ( .A(n6946), .Q(n6945) );
  AOI220 U4590 ( .A(n6329), .B(data_2[6]), .C(n5815), .D(ram_adr[6]), .Q(n4431) );
  NAND30 U4591 ( .A(n1986), .B(n5734), .C(n5699), .Q(n6241) );
  INV3 U4592 ( .A(n6241), .Q(n6242) );
  CLKIN1 U4593 ( .A(n3752), .Q(n1278) );
  AOI221 U4594 ( .A(n1323), .B(n3892), .C(n3866), .D(n3720), .Q(n3891) );
  AOI220 U4595 ( .A(n6509), .B(n1461), .C(n6506), .D(n1460), .Q(n4354) );
  OAI220 U4596 ( .A(n3569), .B(n6258), .C(n1277), .D(n3570), .Q(n4089) );
  INV1 U4597 ( .A(n3863), .Q(n1323) );
  OAI222 U4598 ( .A(n1385), .B(n3973), .C(n3974), .D(n3975), .Q(n3914) );
  CLKIN2 U4599 ( .A(n3983), .Q(n1217) );
  OAI210 U4600 ( .A(n4458), .B(n1310), .C(n4401), .Q(
        \execute/alu/sll_175/temp_int_SH[1] ) );
  NOR21 U4601 ( .A(n3851), .B(n3850), .Q(n3846) );
  MAJ31 U4602 ( .A(n4284), .B(n4285), .C(n4286), .Q(n4283) );
  AOI211 U4603 ( .A(n5696), .B(n4407), .C(n4408), .Q(n4406) );
  INV3 U4604 ( .A(n1772), .Q(n1149) );
  INV6 U4605 ( .A(n6251), .Q(n6252) );
  XNR22 U4606 ( .A(write_register_ex[3]), .B(n1489), .Q(n4570) );
  NOR40 U4607 ( .A(n1771), .B(n1772), .C(n5730), .D(n5716), .Q(n1770) );
  NOR31 U4608 ( .A(n1772), .B(n5730), .C(n6086), .Q(n1773) );
  NAND31 U4609 ( .A(n6246), .B(n6247), .C(n5697), .Q(n6245) );
  OAI2111 U4610 ( .A(n5696), .B(n4417), .C(n4418), .D(n5695), .Q(n4408) );
  OAI211 U4611 ( .A(n4419), .B(n4417), .C(n5946), .Q(n4418) );
  NAND22 U4612 ( .A(n6762), .B(n5731), .Q(n6248) );
  INV3 U4613 ( .A(n6248), .Q(n6249) );
  BUF6 U4614 ( .A(n3475), .Q(n6250) );
  NAND24 U4615 ( .A(n1317), .B(n6236), .Q(n3445) );
  INV6 U4616 ( .A(n6278), .Q(n6312) );
  INV2 U4617 ( .A(n3816), .Q(n1267) );
  AOI220 U4618 ( .A(n1293), .B(n1457), .C(n1289), .D(n1458), .Q(n4353) );
  CLKIN3 U4619 ( .A(n3636), .Q(n1380) );
  AOI220 U4620 ( .A(n6510), .B(n1450), .C(n6506), .D(n1449), .Q(n4193) );
  CLKIN1 U4621 ( .A(n3660), .Q(n1307) );
  CLKIN6 U4622 ( .A(n4543), .Q(n1492) );
  INV2 U4623 ( .A(n4176), .Q(n1366) );
  CLKIN3 U4624 ( .A(n3491), .Q(n1236) );
  INV0 U4625 ( .A(n4170), .Q(n1367) );
  CLKIN6 U4626 ( .A(n6938), .Q(n6936) );
  INV2 U4627 ( .A(n6295), .Q(n6299) );
  AOI221 U4628 ( .A(n1839), .B(pc_out[2]), .C(n1840), .D(inst_out[0]), .Q(
        n1838) );
  AOI221 U4629 ( .A(n6503), .B(write_data_reg[26]), .C(pc_ex[26]), .D(n6323), 
        .Q(n4507) );
  AOI221 U4630 ( .A(n6504), .B(write_data_reg[14]), .C(pc_ex[14]), .D(n6324), 
        .Q(n4492) );
  AOI220 U4631 ( .A(n1467), .B(n6072), .C(pc_ex[1]), .D(n6323), .Q(n4468) );
  AOI220 U4632 ( .A(n6330), .B(data_2[17]), .C(n5816), .D(ram_adr[17]), .Q(
        n4450) );
  NOR42 U4633 ( .A(n2857), .B(n2858), .C(n2859), .D(n2860), .Q(n2856) );
  NOR20 U4634 ( .A(n1459), .B(n6490), .Q(n4285) );
  AOI221 U4635 ( .A(ram_adr[30]), .B(n6336), .C(n6339), .D(data_1[30]), .Q(
        n4528) );
  AOI221 U4636 ( .A(ram_adr[27]), .B(n6336), .C(n6339), .D(data_1[27]), .Q(
        n4523) );
  CLKIN2 U4637 ( .A(n6314), .Q(n6292) );
  INV3 U4638 ( .A(n6290), .Q(n6293) );
  INV3 U4639 ( .A(n6295), .Q(n6298) );
  OAI221 U4640 ( .A(n1243), .B(n3431), .C(n1281), .D(n3554), .Q(n4185) );
  INV2 U4641 ( .A(\execute/alu/sll_175/ML_int[2][0] ), .Q(n1214) );
  OAI222 U4642 ( .A(n1266), .B(n3416), .C(n1267), .D(n3417), .Q(n3450) );
  IMUX20 U4643 ( .A(n6257), .B(n4381), .S(n6343), .Q(
        \execute/alu/sll_175/ML_int[5][16] ) );
  NAND20 U4644 ( .A(n5808), .B(n6756), .Q(n4381) );
  CLKIN2 U4645 ( .A(n3948), .Q(n1225) );
  NOR21 U4646 ( .A(n3569), .B(n5819), .Q(n3507) );
  AOI210 U4647 ( .A(n4058), .B(n1299), .C(n4061), .Q(n4080) );
  AOI220 U4648 ( .A(n6355), .B(n1453), .C(n1294), .D(n1451), .Q(n4249) );
  AOI220 U4649 ( .A(n6353), .B(n1461), .C(n1294), .D(n1458), .Q(n4392) );
  INV2 U4650 ( .A(n5812), .Q(n1216) );
  AOI220 U4651 ( .A(n6355), .B(n1458), .C(n1294), .D(n1456), .Q(n4254) );
  AOI221 U4652 ( .A(n6510), .B(n1460), .C(n6507), .D(n1458), .Q(n4202) );
  AOI220 U4653 ( .A(n6353), .B(n1457), .C(n1294), .D(n1454), .Q(n4146) );
  AOI220 U4654 ( .A(n6355), .B(n1448), .C(n1294), .D(n1445), .Q(n4152) );
  AOI220 U4655 ( .A(n6353), .B(n1447), .C(n1294), .D(n1443), .Q(n4386) );
  AOI220 U4656 ( .A(n6355), .B(n1428), .C(n1294), .D(n1426), .Q(n3606) );
  AOI220 U4657 ( .A(n6355), .B(n1454), .C(n1294), .D(n1452), .Q(n4187) );
  AOI220 U4658 ( .A(n6355), .B(n1426), .C(n1294), .D(n6193), .Q(n3941) );
  CLKIN3 U4659 ( .A(n4019), .Q(n1303) );
  NOR22 U4660 ( .A(n1429), .B(n1366), .Q(n4172) );
  OAI2111 U4661 ( .A(n1406), .B(n3739), .C(n3740), .D(n3741), .Q(n3738) );
  NAND22 U4662 ( .A(n1344), .B(n4366), .Q(n6255) );
  INV3 U4663 ( .A(n6255), .Q(n6256) );
  INV2 U4664 ( .A(n6068), .Q(n6923) );
  NOR24 U4665 ( .A(n1869), .B(n1870), .Q(n1868) );
  INV2 U4666 ( .A(n3622), .Q(n1461) );
  NOR21 U4667 ( .A(n1290), .B(n5821), .Q(n3616) );
  AOI221 U4668 ( .A(n6193), .B(n6512), .C(n3496), .D(n1321), .Q(n3495) );
  AOI220 U4669 ( .A(n1325), .B(n3482), .C(n1349), .D(n3612), .Q(n3576) );
  INV2 U4670 ( .A(n4091), .Q(n1378) );
  NAND20 U4671 ( .A(n3435), .B(n1426), .Q(n3434) );
  OAI210 U4672 ( .A(n3695), .B(n3596), .C(n3696), .Q(n3694) );
  OAI220 U4673 ( .A(n3759), .B(n3390), .C(n1277), .D(n3534), .Q(n4203) );
  AOI220 U4674 ( .A(n6353), .B(n1452), .C(n1294), .D(n1450), .Q(n4148) );
  INV2 U4675 ( .A(n4226), .Q(n1295) );
  AOI220 U4676 ( .A(n6355), .B(n1451), .C(n1294), .D(n1449), .Q(n4390) );
  AOI220 U4677 ( .A(n6510), .B(n1452), .C(n6507), .D(n1451), .Q(n4124) );
  AOI220 U4678 ( .A(n6353), .B(n1449), .C(n1294), .D(n1447), .Q(n4228) );
  AOI220 U4679 ( .A(n6509), .B(n1451), .C(n6506), .D(n1450), .Q(n4359) );
  AOI221 U4680 ( .A(n1315), .B(n3423), .C(\execute/alu/sll_175/ML_int[4][9] ), 
        .D(n1341), .Q(n3422) );
  INV2 U4681 ( .A(n3516), .Q(n1302) );
  NAND22 U4682 ( .A(n5734), .B(\execute/op_21 [17]), .Q(n4018) );
  NAND22 U4683 ( .A(n5734), .B(\execute/op_21 [18]), .Q(n3999) );
  INV2 U4684 ( .A(n4339), .Q(n1384) );
  NAND22 U4685 ( .A(n5734), .B(\execute/op_21 [20]), .Q(n3911) );
  NAND22 U4686 ( .A(n5734), .B(\execute/op_21 [19]), .Q(n3972) );
  AOI222 U4687 ( .A(n6072), .B(n6490), .C(\execute/op_21 [7]), .D(n5734), .Q(
        n3465) );
  INV2 U4688 ( .A(n4338), .Q(n1370) );
  AOI2110 U4689 ( .A(n3402), .B(n5817), .C(n3684), .D(n6512), .Q(n3682) );
  AOI210 U4690 ( .A(n6512), .B(n5817), .C(n3694), .Q(n3677) );
  AOI220 U4691 ( .A(\execute/alu/sll_175/ML_int[5][20] ), .B(n1353), .C(n6236), 
        .D(n3572), .Q(n3900) );
  CLKIN0 U4692 ( .A(n6341), .Q(n1259) );
  NOR40 U4693 ( .A(n3411), .B(n3412), .C(n1339), .D(n3413), .Q(n3409) );
  XNR20 U4694 ( .A(n3418), .B(n1297), .Q(n3408) );
  AOI220 U4695 ( .A(n6355), .B(n6222), .C(n1294), .D(n5830), .Q(n4142) );
  AOI220 U4696 ( .A(n6355), .B(n5829), .C(n1294), .D(n6346), .Q(n4373) );
  AOI220 U4697 ( .A(n6353), .B(n6346), .C(n1294), .D(n6344), .Q(n4257) );
  AOI220 U4698 ( .A(n6355), .B(n6345), .C(n1294), .D(n1428), .Q(n3946) );
  AOI220 U4699 ( .A(\execute/alu/sll_175/ML_int[5][19] ), .B(n1353), .C(n6236), 
        .D(n3612), .Q(n3960) );
  AOI220 U4700 ( .A(n6355), .B(n6344), .C(n1294), .D(n1427), .Q(n4378) );
  AOI220 U4701 ( .A(n6356), .B(n6346), .C(n1294), .D(n6345), .Q(n4206) );
  OAI220 U4702 ( .A(n3595), .B(n3596), .C(n3569), .D(n1855), .Q(n3594) );
  AOI220 U4703 ( .A(n6355), .B(n1443), .C(n1294), .D(n5829), .Q(n4252) );
  AOI220 U4704 ( .A(n6510), .B(n6345), .C(n6507), .D(n6344), .Q(n3956) );
  AOI220 U4705 ( .A(n3602), .B(n1443), .C(n1294), .D(n6222), .Q(n4191) );
  AOI220 U4706 ( .A(n6329), .B(data_2[7]), .C(n5815), .D(ram_adr[7]), .Q(n4430) );
  BUF15 U4707 ( .A(\execute/n432 ), .Q(n6346) );
  INV4 U4708 ( .A(\execute/op_21 [13]), .Q(n1435) );
  OAI222 U4709 ( .A(n5107), .B(n6566), .C(n5106), .D(n6563), .Q(n3179) );
  OAI222 U4710 ( .A(n5301), .B(n6567), .C(n5300), .D(n6563), .Q(n3137) );
  OAI222 U4711 ( .A(n5299), .B(n6576), .C(n5298), .D(n1928), .Q(n3138) );
  OAI222 U4712 ( .A(n5109), .B(n6557), .C(n5108), .D(n6554), .Q(n3178) );
  OAI222 U4713 ( .A(n5303), .B(n6558), .C(n5302), .D(n6554), .Q(n3136) );
  OAI222 U4714 ( .A(n5255), .B(n6535), .C(n5254), .D(n6528), .Q(n2049) );
  OAI222 U4715 ( .A(n5147), .B(n6529), .C(n5146), .D(n6527), .Q(n2658) );
  OAI222 U4716 ( .A(n5169), .B(n6530), .C(n5168), .D(n6528), .Q(n2511) );
  OAI222 U4717 ( .A(n5145), .B(n6538), .C(n5144), .D(n6537), .Q(n2659) );
  OAI222 U4718 ( .A(n5171), .B(n6521), .C(n5170), .D(n6519), .Q(n2510) );
  OAI222 U4719 ( .A(n5227), .B(n6521), .C(n5226), .D(n6519), .Q(n2531) );
  INV3 U4720 ( .A(write_data_reg[27]), .Q(n6986) );
  AOI220 U4721 ( .A(n6330), .B(data_2[9]), .C(n5815), .D(ram_adr[9]), .Q(n4426) );
  INV3 U4722 ( .A(write_data_reg[18]), .Q(n6968) );
  OAI222 U4723 ( .A(n4953), .B(n6578), .C(n4952), .D(n1928), .Q(n2890) );
  AOI2111 U4724 ( .A(n5544), .B(n6389), .C(n2872), .D(n2873), .Q(n2855) );
  AOI2111 U4725 ( .A(n5520), .B(n6386), .C(n2935), .D(n2936), .Q(n2918) );
  AOI2111 U4726 ( .A(n5512), .B(n6391), .C(n2956), .D(n2957), .Q(n2939) );
  AOI2111 U4727 ( .A(n5496), .B(n6391), .C(n2998), .D(n2999), .Q(n2981) );
  AOI221 U4728 ( .A(n6364), .B(n5908), .C(n5494), .D(n1954), .Q(n2979) );
  AOI2111 U4729 ( .A(n5536), .B(n6452), .C(n2204), .D(n2205), .Q(n2187) );
  OAI222 U4730 ( .A(n4891), .B(n6585), .C(n4890), .D(n6582), .Q(n3181) );
  OAI222 U4731 ( .A(n5305), .B(n6586), .C(n5304), .D(n6582), .Q(n3139) );
  AOI2111 U4732 ( .A(n5528), .B(n6387), .C(n2914), .D(n2915), .Q(n2897) );
  AOI2111 U4733 ( .A(n5536), .B(n6388), .C(n2893), .D(n2894), .Q(n2876) );
  OAI222 U4734 ( .A(n5105), .B(n6575), .C(n5104), .D(n6573), .Q(n3180) );
  OAI222 U4735 ( .A(n4905), .B(n6547), .C(n4904), .D(n6545), .Q(n2660) );
  OAI222 U4736 ( .A(n4977), .B(n6575), .C(n4976), .D(n6572), .Q(n3184) );
  OAI222 U4737 ( .A(n5295), .B(n6567), .C(n5294), .D(n6563), .Q(n3141) );
  OAI222 U4738 ( .A(n5293), .B(n6576), .C(n5292), .D(n1928), .Q(n3142) );
  OAI222 U4739 ( .A(n4877), .B(n6551), .C(n4876), .D(n2009), .Q(n2303) );
  OAI222 U4740 ( .A(n4885), .B(n6548), .C(n4884), .D(n6545), .Q(n2576) );
  OAI222 U4741 ( .A(n4923), .B(n6547), .C(n4922), .D(n6545), .Q(n2618) );
  OAI222 U4742 ( .A(n4937), .B(n6547), .C(n4936), .D(n6545), .Q(n2639) );
  OAI222 U4743 ( .A(n5003), .B(n6571), .C(n5002), .D(n6564), .Q(n1934) );
  OAI222 U4744 ( .A(n5001), .B(n6580), .C(n5000), .D(n1928), .Q(n1935) );
  OAI222 U4745 ( .A(n4913), .B(n6548), .C(n4912), .D(n2009), .Q(n2513) );
  OAI222 U4746 ( .A(n4929), .B(n6548), .C(n4928), .D(n6545), .Q(n2534) );
  OAI222 U4747 ( .A(n4939), .B(n6553), .C(n4938), .D(n6546), .Q(n2051) );
  OAI222 U4748 ( .A(n5297), .B(n6558), .C(n5296), .D(n6554), .Q(n3140) );
  OAI222 U4749 ( .A(n5005), .B(n6562), .C(n5004), .D(n6555), .Q(n1933) );
  OAI222 U4750 ( .A(n5253), .B(n6544), .C(n5252), .D(n6537), .Q(n2050) );
  OAI222 U4751 ( .A(n5125), .B(n6535), .C(n5124), .D(n2013), .Q(n2053) );
  OAI222 U4752 ( .A(n5123), .B(n6544), .C(n5122), .D(n6537), .Q(n2054) );
  OAI222 U4753 ( .A(n5059), .B(n6533), .C(n5058), .D(n6527), .Q(n2301) );
  OAI222 U4754 ( .A(n5057), .B(n6542), .C(n5056), .D(n6536), .Q(n2302) );
  OAI222 U4755 ( .A(n4965), .B(n6542), .C(n4964), .D(n6537), .Q(n2306) );
  OAI222 U4756 ( .A(n5225), .B(n6530), .C(n5224), .D(n6528), .Q(n2532) );
  OAI222 U4757 ( .A(n5167), .B(n6539), .C(n5166), .D(n6536), .Q(n2512) );
  OAI222 U4758 ( .A(n5223), .B(n6539), .C(n5222), .D(n6536), .Q(n2533) );
  OAI222 U4759 ( .A(n4999), .B(n6529), .C(n4998), .D(n6527), .Q(n2662) );
  OAI222 U4760 ( .A(n5083), .B(n6530), .C(n5082), .D(n6527), .Q(n2574) );
  OAI222 U4761 ( .A(n4997), .B(n6538), .C(n4996), .D(n2011), .Q(n2663) );
  OAI222 U4762 ( .A(n5081), .B(n6539), .C(n5080), .D(n6536), .Q(n2575) );
  OAI222 U4763 ( .A(n5071), .B(n6530), .C(n5070), .D(n6528), .Q(n2536) );
  OAI222 U4764 ( .A(n5011), .B(n6539), .C(n5010), .D(n6536), .Q(n2516) );
  OAI222 U4765 ( .A(n5209), .B(n6529), .C(n5208), .D(n6527), .Q(n2616) );
  OAI222 U4766 ( .A(n5069), .B(n6539), .C(n5068), .D(n6536), .Q(n2537) );
  OAI222 U4767 ( .A(n5207), .B(n6538), .C(n5206), .D(n2011), .Q(n2617) );
  OAI222 U4768 ( .A(n5249), .B(n6529), .C(n5248), .D(n6527), .Q(n2637) );
  OAI222 U4769 ( .A(n4971), .B(n6530), .C(n4970), .D(n6527), .Q(n2578) );
  OAI222 U4770 ( .A(n5247), .B(n6538), .C(n5246), .D(n2011), .Q(n2638) );
  OAI222 U4771 ( .A(n4969), .B(n6539), .C(n4968), .D(n6536), .Q(n2579) );
  OAI222 U4772 ( .A(n5053), .B(n6529), .C(n5052), .D(n6527), .Q(n2620) );
  OAI222 U4773 ( .A(n5051), .B(n6538), .C(n5050), .D(n2011), .Q(n2621) );
  OAI222 U4774 ( .A(n5113), .B(n6529), .C(n5112), .D(n6527), .Q(n2641) );
  OAI222 U4775 ( .A(n5111), .B(n6538), .C(n5110), .D(n2011), .Q(n2642) );
  OAI222 U4776 ( .A(n5339), .B(n6524), .C(n5338), .D(n2015), .Q(n2304) );
  OAI222 U4777 ( .A(n5085), .B(n6521), .C(n5084), .D(n6518), .Q(n2573) );
  OAI222 U4778 ( .A(n5015), .B(n6521), .C(n5014), .D(n6519), .Q(n2514) );
  OAI222 U4779 ( .A(n5073), .B(n6521), .C(n5072), .D(n6519), .Q(n2535) );
  OAI222 U4780 ( .A(n5211), .B(n6520), .C(n5210), .D(n6518), .Q(n2615) );
  OAI222 U4781 ( .A(n5251), .B(n6520), .C(n5250), .D(n6518), .Q(n2636) );
  OAI222 U4782 ( .A(n5313), .B(n6521), .C(n5312), .D(n6518), .Q(n2577) );
  OAI222 U4783 ( .A(n5055), .B(n6520), .C(n5054), .D(n6518), .Q(n2619) );
  OAI222 U4784 ( .A(n5115), .B(n6520), .C(n5114), .D(n6518), .Q(n2640) );
  OAI220 U4785 ( .A(n4659), .B(n6414), .C(n4658), .D(n6416), .Q(n2900) );
  OAI220 U4786 ( .A(n4583), .B(n1939), .C(n4582), .D(n1940), .Q(n2858) );
  OAI220 U4787 ( .A(n4603), .B(n1939), .C(n4602), .D(n1940), .Q(n2984) );
  NOR41 U4788 ( .A(n2863), .B(n2864), .C(n2865), .D(n2866), .Q(n2862) );
  INV0 U4789 ( .A(n3445), .Q(n1315) );
  OAI220 U4790 ( .A(n1267), .B(n3570), .C(n1227), .D(n3445), .Q(n3731) );
  IMUX20 U4791 ( .A(\execute/alu/sll_175/ML_int[3][15] ), .B(
        \execute/alu/sll_175/ML_int[3][7] ), .S(n5819), .Q(n6258) );
  CLKIN3 U4792 ( .A(n6511), .Q(n6510) );
  CLKIN3 U4793 ( .A(n6508), .Q(n6506) );
  CLKIN2 U4794 ( .A(n6508), .Q(n6507) );
  AOI310 U4795 ( .A(n1341), .B(n5819), .C(\execute/alu/sll_175/ML_int[3][14] ), 
        .D(n1348), .Q(n3881) );
  IMUX20 U4796 ( .A(\execute/alu/sll_175/ML_int[3][16] ), .B(
        \execute/alu/sll_175/ML_int[3][8] ), .S(n5819), .Q(n6257) );
  INV0 U4797 ( .A(n3775), .Q(n1274) );
  OAI220 U4798 ( .A(n1230), .B(n3430), .C(n1231), .D(n3431), .Q(n3429) );
  OAI220 U4799 ( .A(n1280), .B(n3416), .C(n1278), .D(n3417), .Q(n3479) );
  OAI220 U4800 ( .A(n1245), .B(n3431), .C(n1280), .D(n3554), .Q(n4075) );
  OAI220 U4801 ( .A(n1286), .B(n3416), .C(n1288), .D(n3417), .Q(n3411) );
  NAND20 U4802 ( .A(n5810), .B(n6759), .Q(n3948) );
  IMUX20 U4803 ( .A(n6259), .B(n1856), .S(n6343), .Q(
        \execute/alu/sll_175/ML_int[5][20] ) );
  IMUX20 U4804 ( .A(n6260), .B(n1855), .S(n6343), .Q(
        \execute/alu/sll_175/ML_int[5][19] ) );
  INV0 U4805 ( .A(n3454), .Q(n1322) );
  CLKIN3 U4806 ( .A(n3487), .Q(n1211) );
  NAND20 U4807 ( .A(n3673), .B(n1306), .Q(n3743) );
  CLKIN3 U4808 ( .A(n3529), .Q(n1221) );
  INV0 U4809 ( .A(n3624), .Q(n1254) );
  CLKIN6 U4810 ( .A(n6505), .Q(n6503) );
  INV0 U4811 ( .A(n3641), .Q(n1400) );
  AOI210 U4812 ( .A(n4139), .B(n4140), .C(n4059), .Q(n4129) );
  INV1 U4813 ( .A(n3867), .Q(n1270) );
  NAND20 U4814 ( .A(n1349), .B(n1317), .Q(n4082) );
  OAI210 U4815 ( .A(n3667), .B(n3633), .C(n3643), .Q(n3660) );
  AOI220 U4816 ( .A(n1293), .B(n1450), .C(n1289), .D(n1451), .Q(n4273) );
  AOI220 U4817 ( .A(n6509), .B(n1453), .C(n6506), .D(n1452), .Q(n4274) );
  AOI220 U4818 ( .A(n1293), .B(n1456), .C(n1289), .D(n1457), .Q(n4201) );
  AOI220 U4819 ( .A(n1313), .B(n3395), .C(n1333), .D(n3800), .Q(n4114) );
  AOI220 U4820 ( .A(n1335), .B(n3396), .C(n1325), .D(n3544), .Q(n4113) );
  AOI2110 U4821 ( .A(\execute/alu/sll_175/ML_int[4][13] ), .B(n1341), .C(n4141), .D(n4102), .Q(n4115) );
  AOI220 U4822 ( .A(n1313), .B(n3921), .C(n1333), .D(n3815), .Q(n4155) );
  AOI220 U4823 ( .A(n1335), .B(n3575), .C(n1325), .D(n3557), .Q(n4154) );
  AOI2110 U4824 ( .A(\execute/alu/sll_175/ML_int[4][12] ), .B(n1341), .C(n4177), .D(n4102), .Q(n4156) );
  AOI220 U4825 ( .A(n1313), .B(n3862), .C(n1333), .D(n3861), .Q(n4093) );
  AOI220 U4826 ( .A(n1331), .B(n3775), .C(n1328), .D(n3867), .Q(n4094) );
  NOR30 U4827 ( .A(n1342), .B(n5819), .C(n4006), .Q(n3878) );
  NAND20 U4828 ( .A(n3802), .B(n3899), .Q(n3871) );
  OAI210 U4829 ( .A(n3739), .B(n1306), .C(n3764), .Q(n3778) );
  NAND20 U4830 ( .A(n3805), .B(n3802), .Q(n3826) );
  INV0 U4831 ( .A(n4401), .Q(n1359) );
  AOI220 U4832 ( .A(n4169), .B(n1298), .C(n1369), .D(n4140), .Q(n4167) );
  NOR20 U4833 ( .A(n1369), .B(n4059), .Q(n4169) );
  AOI220 U4834 ( .A(n1293), .B(n1453), .C(n1289), .D(n1454), .Q(n4121) );
  AOI220 U4835 ( .A(n1293), .B(n6222), .C(n1289), .D(n1443), .Q(n4360) );
  AOI220 U4836 ( .A(n6509), .B(n1447), .C(n6506), .D(n1445), .Q(n4361) );
  AOI220 U4837 ( .A(n1293), .B(n1452), .C(n1289), .D(n1453), .Q(n4356) );
  AOI220 U4838 ( .A(n6509), .B(n1456), .C(n6506), .D(n1454), .Q(n4357) );
  AOI220 U4839 ( .A(n1293), .B(n1443), .C(n1289), .D(n1445), .Q(n4150) );
  AOI220 U4840 ( .A(n6510), .B(n1448), .C(n6506), .D(n1447), .Q(n4151) );
  AOI220 U4841 ( .A(n4138), .B(n4129), .C(n1371), .D(n1299), .Q(n4136) );
  NOR20 U4842 ( .A(n1371), .B(n4061), .Q(n4138) );
  NAND20 U4843 ( .A(n3834), .B(n1330), .Q(n3864) );
  NOR20 U4844 ( .A(n1242), .B(n3445), .Q(n4204) );
  NAND20 U4845 ( .A(n1461), .B(n3863), .Q(n3765) );
  OAI220 U4846 ( .A(n1268), .B(n3570), .C(n1234), .D(n3445), .Q(n4177) );
  OAI220 U4847 ( .A(n1272), .B(n3570), .C(n1237), .D(n3445), .Q(n4099) );
  NAND20 U4848 ( .A(n1386), .B(n3912), .Q(n3969) );
  XNR20 U4849 ( .A(n3802), .B(n3909), .Q(n3908) );
  NOR20 U4850 ( .A(n1390), .B(n3872), .Q(n3909) );
  OAI212 U4851 ( .A(n3773), .B(n3596), .C(n3774), .Q(n3771) );
  AOI220 U4852 ( .A(n1323), .B(n3557), .C(n1327), .D(n3917), .Q(n4351) );
  AOI220 U4853 ( .A(n3866), .B(n3817), .C(n3994), .D(n3816), .Q(n4352) );
  AOI220 U4854 ( .A(n1349), .B(n3486), .C(n1211), .D(n1341), .Q(n3456) );
  INV0 U4855 ( .A(n4140), .Q(n1298) );
  INV0 U4856 ( .A(n3513), .Q(n1271) );
  XNR20 U4857 ( .A(n3801), .B(n3667), .Q(n3799) );
  OAI222 U4858 ( .A(n3407), .B(n3799), .C(n3391), .D(n3596), .Q(n3798) );
  OAI220 U4859 ( .A(n1269), .B(n3534), .C(n1232), .D(n3535), .Q(n3566) );
  OAI220 U4860 ( .A(n1231), .B(n3430), .C(n1234), .D(n3431), .Q(n3565) );
  NOR20 U4861 ( .A(n1305), .B(n3725), .Q(n3736) );
  OAI221 U4862 ( .A(n1265), .B(n3553), .C(n1268), .D(n3554), .Q(n3552) );
  AOI220 U4863 ( .A(n1293), .B(n1451), .C(n1289), .D(n1452), .Q(n4198) );
  AOI220 U4864 ( .A(n6510), .B(n1454), .C(n6506), .D(n1453), .Q(n4199) );
  AOI220 U4865 ( .A(n1292), .B(n3994), .C(n3866), .D(n3775), .Q(n3992) );
  OAI220 U4866 ( .A(n1283), .B(n3415), .C(n1287), .D(n1322), .Q(n3412) );
  OAI210 U4867 ( .A(n1394), .B(n3871), .C(n3848), .Q(n3868) );
  INV0 U4868 ( .A(n3640), .Q(n1397) );
  AOI220 U4869 ( .A(n1323), .B(n3544), .C(n3866), .D(n3797), .Q(n4027) );
  AOI220 U4870 ( .A(n1327), .B(n3892), .C(n3994), .D(n3720), .Q(n4026) );
  AOI220 U4871 ( .A(n1293), .B(n1425), .C(n1289), .D(n1426), .Q(n3613) );
  AOI220 U4872 ( .A(n3615), .B(n1428), .C(n6507), .D(n1427), .Q(n3614) );
  AOI220 U4873 ( .A(n1293), .B(n1422), .C(n1289), .D(n6193), .Q(n3957) );
  AOI220 U4874 ( .A(n3615), .B(n1426), .C(n6507), .D(n1425), .Q(n3958) );
  AOI220 U4875 ( .A(n1293), .B(n6193), .C(n1289), .D(n1425), .Q(n3707) );
  AOI220 U4876 ( .A(n3615), .B(n1427), .C(n6507), .D(n1426), .Q(n3708) );
  INV0 U4877 ( .A(n3485), .Q(n1281) );
  CLKIN1 U4878 ( .A(n3917), .Q(n1264) );
  INV0 U4879 ( .A(n3872), .Q(n1391) );
  CLKIN3 U4880 ( .A(n4463), .Q(n1224) );
  NAND20 U4881 ( .A(\execute/alu/sll_175/ML_int[2][3] ), .B(n6759), .Q(n4463)
         );
  INV2 U4882 ( .A(n4092), .Q(n1241) );
  AOI220 U4883 ( .A(n3814), .B(n1336), .C(n3815), .D(n1317), .Q(n3446) );
  AOI220 U4884 ( .A(n6356), .B(n1452), .C(n1450), .D(n1258), .Q(n4250) );
  AOI220 U4885 ( .A(n6356), .B(n1460), .C(n1457), .D(n1258), .Q(n4393) );
  AOI220 U4886 ( .A(n6356), .B(n1457), .C(n1454), .D(n1258), .Q(n4255) );
  AOI220 U4887 ( .A(n3602), .B(n1454), .C(n1452), .D(n1258), .Q(n4389) );
  AOI220 U4888 ( .A(n3602), .B(n1456), .C(n1453), .D(n1258), .Q(n4147) );
  AOI220 U4889 ( .A(n6356), .B(n1445), .C(n6222), .D(n1258), .Q(n4387) );
  AOI220 U4890 ( .A(n1317), .B(n3396), .C(n1334), .D(n3713), .Q(n4028) );
  NAND20 U4891 ( .A(n3639), .B(n3640), .Q(n3804) );
  AOI220 U4892 ( .A(n6356), .B(n1453), .C(n1451), .D(n1258), .Q(n4188) );
  AOI220 U4893 ( .A(n1317), .B(n3501), .C(n1336), .D(n3862), .Q(n3990) );
  AOI220 U4894 ( .A(n1314), .B(n3815), .C(n1317), .D(n3575), .Q(n4385) );
  AOI220 U4895 ( .A(n3602), .B(n1425), .C(n1258), .D(n1422), .Q(n3942) );
  AOI220 U4896 ( .A(n3664), .B(n1336), .C(n3861), .D(n1317), .Q(n3773) );
  AOI220 U4897 ( .A(n3837), .B(n1317), .C(n1254), .D(n1336), .Q(n3759) );
  AOI220 U4898 ( .A(n3713), .B(n1336), .C(n3800), .D(n1317), .Q(n3391) );
  AOI220 U4899 ( .A(n3602), .B(n1447), .C(n1443), .D(n1258), .Q(n4153) );
  AOI220 U4900 ( .A(n6356), .B(n1427), .C(n1258), .D(n1425), .Q(n3607) );
  AOI220 U4901 ( .A(n6355), .B(n1427), .C(n1294), .D(n1425), .Q(n3703) );
  AOI220 U4902 ( .A(n6356), .B(n1426), .C(n1258), .D(n6193), .Q(n3704) );
  AOI220 U4903 ( .A(n1317), .B(n3981), .C(n1336), .D(n3982), .Q(n3979) );
  INV0 U4904 ( .A(n3642), .Q(n1399) );
  INV0 U4905 ( .A(n3671), .Q(n1403) );
  INV2 U4906 ( .A(n6068), .Q(n6924) );
  CLKIN3 U4907 ( .A(n1985), .Q(n1145) );
  NOR20 U4908 ( .A(n6261), .B(n1377), .Q(n4047) );
  XNR20 U4909 ( .A(n3745), .B(n6350), .Q(n3726) );
  XNR20 U4910 ( .A(n3659), .B(n6321), .Q(n3662) );
  XNR20 U4911 ( .A(n3999), .B(n6351), .Q(n3973) );
  NOR20 U4912 ( .A(n4020), .B(n1383), .Q(n4001) );
  XNR20 U4913 ( .A(n3781), .B(n3627), .Q(n3786) );
  XNR20 U4914 ( .A(n3972), .B(n6350), .Q(n3970) );
  XNR20 U4915 ( .A(n3821), .B(n6351), .Q(n3825) );
  NAND20 U4916 ( .A(n3806), .B(n1404), .Q(n3764) );
  CLKIN6 U4917 ( .A(n3587), .Q(n1417) );
  INV0 U4918 ( .A(n4055), .Q(n1350) );
  AOI210 U4919 ( .A(n3515), .B(n3516), .C(n3517), .Q(n3474) );
  NOR20 U4920 ( .A(n3622), .B(n4270), .Q(n3834) );
  CLKIN1 U4921 ( .A(n3538), .Q(n1422) );
  AOI220 U4922 ( .A(n1293), .B(n1458), .C(n1289), .D(n1460), .Q(n4135) );
  AOI220 U4923 ( .A(n3497), .B(n1315), .C(n3498), .D(n1349), .Q(n3494) );
  AOI220 U4924 ( .A(n3499), .B(n1325), .C(n3500), .D(n1335), .Q(n3493) );
  AOI220 U4925 ( .A(n3646), .B(n6352), .C(n6358), .D(n3622), .Q(n3645) );
  OAI2110 U4926 ( .A(n1439), .B(n3617), .C(n3618), .D(n3619), .Q(
        \execute/old_res [31]) );
  NOR20 U4927 ( .A(n3561), .B(n1352), .Q(n3527) );
  NAND21 U4928 ( .A(n4270), .B(n1330), .Q(n3890) );
  NAND30 U4929 ( .A(n1383), .B(n4018), .C(n1470), .Q(n4022) );
  AOI220 U4930 ( .A(n4023), .B(n1303), .C(n1382), .D(n4019), .Q(n4021) );
  NOR20 U4931 ( .A(n1382), .B(n4001), .Q(n4023) );
  OAI2110 U4932 ( .A(n1374), .B(n6352), .C(n1324), .D(n4100), .Q(n4097) );
  AOI220 U4933 ( .A(n1328), .B(n3545), .C(n1347), .D(n3546), .Q(n3521) );
  AOI220 U4934 ( .A(n1313), .B(n3394), .C(n1333), .D(n3396), .Q(n3520) );
  AOI220 U4935 ( .A(n1293), .B(n1445), .C(n1289), .D(n1447), .Q(n4271) );
  AOI220 U4936 ( .A(n6509), .B(n1449), .C(n6506), .D(n1448), .Q(n4272) );
  AOI2110 U4937 ( .A(n1347), .B(n3580), .C(n3581), .D(n3582), .Q(n3579) );
  AOI210 U4938 ( .A(n1315), .B(n3500), .C(n4251), .Q(n4220) );
  AOI2110 U4939 ( .A(n1333), .B(n3862), .C(n4222), .D(n4223), .Q(n4221) );
  AOI220 U4940 ( .A(n1471), .B(n1414), .C(n6512), .D(n6253), .Q(n4032) );
  AOI2110 U4941 ( .A(n1381), .B(n4034), .C(n4035), .D(n4036), .Q(n4033) );
  AOI220 U4942 ( .A(n6516), .B(n1454), .C(n6515), .D(n3781), .Q(n3780) );
  OAI220 U4943 ( .A(n3773), .B(n3390), .C(n1237), .D(n3535), .Q(n4251) );
  OAI220 U4944 ( .A(n1232), .B(n3445), .C(n3446), .D(n3390), .Q(n3444) );
  AOI220 U4945 ( .A(n1361), .B(n1426), .C(n1360), .D(n1425), .Q(n4337) );
  AOI2110 U4946 ( .A(n1300), .B(n3476), .C(n1219), .D(n3503), .Q(n3490) );
  OAI310 U4947 ( .A(n3407), .B(n3474), .C(n6250), .D(n3504), .Q(n3503) );
  AOI220 U4948 ( .A(n1293), .B(n1449), .C(n1289), .D(n1450), .Q(n4123) );
  AOI220 U4949 ( .A(n1293), .B(n1447), .C(n1289), .D(n1448), .Q(n4192) );
  AOI220 U4950 ( .A(n1293), .B(n1448), .C(n1289), .D(n1449), .Q(n4358) );
  OAI310 U4951 ( .A(n3407), .B(n3474), .C(n3476), .D(n3510), .Q(n3509) );
  AOI220 U4952 ( .A(n3506), .B(n1358), .C(n3507), .D(
        \execute/alu/sll_175/ML_int[3][6] ), .Q(n3505) );
  OAI220 U4953 ( .A(n1244), .B(n3445), .C(n1281), .D(n3534), .Q(n4088) );
  AOI220 U4954 ( .A(n6236), .B(n3931), .C(n1471), .D(n1415), .Q(n4010) );
  AOI2110 U4955 ( .A(n5811), .B(n1341), .C(n3925), .D(n3926), .Q(n3924) );
  OAI210 U4956 ( .A(n4458), .B(n1344), .C(n4401), .Q(
        \execute/alu/sll_175/temp_int_SH[4] ) );
  NOR20 U4957 ( .A(n4047), .B(n1376), .Q(n4078) );
  AOI220 U4958 ( .A(n3394), .B(n1335), .C(n3395), .D(n1333), .Q(n3393) );
  AOI220 U4959 ( .A(\execute/alu/sll_175/ML_int[4][10] ), .B(n1341), .C(n1473), 
        .D(n4259), .Q(n4218) );
  AOI220 U4960 ( .A(n3454), .B(n3499), .C(n3455), .D(n3518), .Q(n4261) );
  AOI220 U4961 ( .A(n1332), .B(n3867), .C(n1329), .D(n3513), .Q(n4260) );
  NAND20 U4962 ( .A(n1319), .B(n3589), .Q(n3688) );
  NAND20 U4963 ( .A(n3635), .B(n1412), .Q(n3661) );
  OAI220 U4964 ( .A(n1243), .B(n3430), .C(n1244), .D(n3431), .Q(n3462) );
  AOI220 U4965 ( .A(n3501), .B(n1333), .C(n3502), .D(n1313), .Q(n3492) );
  OAI220 U4966 ( .A(n1244), .B(n3535), .C(n1245), .D(n3430), .Q(n4186) );
  OAI2110 U4967 ( .A(n1429), .B(n1295), .C(n4230), .D(n4231), .Q(n4222) );
  AOI210 U4968 ( .A(n3701), .B(n3702), .C(n3601), .Q(n3700) );
  OAI2110 U4969 ( .A(n3569), .B(n4381), .C(n4382), .D(n4383), .Q(n4362) );
  NOR20 U4970 ( .A(n3970), .B(n1387), .Q(n3971) );
  AOI220 U4971 ( .A(n1329), .B(n3484), .C(n1332), .D(n3485), .Q(n3483) );
  NAND20 U4972 ( .A(n1392), .B(n3826), .Q(n3845) );
  AOI220 U4973 ( .A(n3481), .B(n3455), .C(n3482), .D(n3454), .Q(n3480) );
  CLKIN2 U4974 ( .A(n3852), .Q(n1220) );
  AOI220 U4975 ( .A(n3954), .B(n1347), .C(n3536), .D(n1328), .Q(n3953) );
  OAI2110 U4976 ( .A(n3745), .B(n4131), .C(n4209), .D(n4210), .Q(n3837) );
  AOI220 U4977 ( .A(n1456), .B(n1258), .C(n3603), .D(n1460), .Q(n4210) );
  NOR20 U4978 ( .A(n4087), .B(n3622), .Q(n4085) );
  AOI220 U4979 ( .A(n3602), .B(n1461), .C(n1458), .D(n1258), .Q(n4132) );
  XOR20 U4980 ( .A(n3440), .B(n3441), .Q(n3432) );
  AOI220 U4981 ( .A(n6356), .B(n1451), .C(n1449), .D(n1258), .Q(n4149) );
  AOI220 U4982 ( .A(n6356), .B(n1450), .C(n1448), .D(n1258), .Q(n4391) );
  AOI310 U4983 ( .A(n6352), .B(n4037), .C(n4038), .D(n1381), .Q(n4036) );
  AOI310 U4984 ( .A(n4016), .B(n6352), .C(n4017), .D(n1383), .Q(n4015) );
  INV0 U4985 ( .A(n4020), .Q(n1444) );
  AOI220 U4986 ( .A(n1317), .B(n3395), .C(n1336), .D(n3800), .Q(n3896) );
  CLKIN1 U4987 ( .A(n3781), .Q(n1454) );
  AOI220 U4988 ( .A(n1447), .B(n1258), .C(n6355), .D(n1450), .Q(n4195) );
  CLKIN1 U4989 ( .A(n3793), .Q(n1453) );
  CLKIN1 U4990 ( .A(n3755), .Q(n1456) );
  CLKIN1 U4991 ( .A(n3843), .Q(n1451) );
  CLKIN1 U4992 ( .A(n3821), .Q(n1452) );
  NOR20 U4993 ( .A(n3622), .B(n6234), .Q(n4086) );
  AOI220 U4994 ( .A(n6356), .B(n1448), .C(n1445), .D(n1258), .Q(n4229) );
  NAND20 U4995 ( .A(n3563), .B(n1351), .Q(n3560) );
  AOI220 U4996 ( .A(n3560), .B(n3561), .C(n3527), .D(n3562), .Q(n3558) );
  NAND30 U4997 ( .A(n1478), .B(n6176), .C(n4064), .Q(n3410) );
  CLKIN1 U4998 ( .A(n3745), .Q(n1457) );
  CLKIN1 U4999 ( .A(n3716), .Q(n1458) );
  CLKIN1 U5000 ( .A(n3870), .Q(n1450) );
  OAI220 U5001 ( .A(n4256), .B(n3659), .C(n3622), .D(n4131), .Q(n3664) );
  CLKIN1 U5002 ( .A(n3659), .Q(n1460) );
  NAND30 U5003 ( .A(n1374), .B(n1436), .C(n1470), .Q(n4106) );
  AOI210 U5004 ( .A(n6515), .B(n1372), .C(n6512), .Q(n4133) );
  NOR20 U5005 ( .A(n3658), .B(n3659), .Q(n3655) );
  OAI210 U5006 ( .A(n1395), .B(n3875), .C(n3874), .Q(n3898) );
  NAND20 U5007 ( .A(n1372), .B(n1434), .Q(n4137) );
  NAND20 U5008 ( .A(n1366), .B(n1429), .Q(n4217) );
  OAI210 U5009 ( .A(n6515), .B(n3622), .C(n1413), .Q(n3646) );
  NOR20 U5010 ( .A(n4350), .B(n4394), .Q(n4367) );
  CLKIN2 U5011 ( .A(n4473), .Q(n1364) );
  CLKBU12 U5012 ( .A(n1841), .Q(n6270) );
  AOI212 U5013 ( .A(n1319), .B(n1417), .C(n1338), .Q(n4245) );
  AOI2112 U5014 ( .A(n3587), .B(n3591), .C(n4245), .D(n4246), .Q(n4054) );
  NAND22 U5015 ( .A(n3562), .B(n3564), .Q(n3563) );
  NAND20 U5016 ( .A(n3850), .B(n3851), .Q(n3849) );
  OAI310 U5017 ( .A(n1187), .B(n1145), .C(n6085), .D(n1146), .Q(
        \instruction_decode/old_wb[1] ) );
  CLKIN1 U5018 ( .A(n3746), .Q(n1409) );
  XOR22 U5019 ( .A(\instruction_decode/old_data_1 [28]), .B(
        \instruction_decode/old_data_2 [28]), .Q(n1909) );
  XOR22 U5020 ( .A(\instruction_decode/old_data_1 [29]), .B(
        \instruction_decode/old_data_2 [29]), .Q(n1908) );
  XOR22 U5021 ( .A(\instruction_decode/old_data_1 [31]), .B(
        \instruction_decode/old_data_2 [31]), .Q(n1888) );
  AOI220 U5022 ( .A(n1453), .B(n1404), .C(n1454), .D(n1405), .Q(n4297) );
  AOI210 U5023 ( .A(n1449), .B(n1395), .C(n4300), .Q(n4304) );
  OAI210 U5024 ( .A(n1422), .B(n1356), .C(n4329), .Q(n4328) );
  XOR22 U5025 ( .A(\instruction_decode/old_data_1 [26]), .B(
        \instruction_decode/old_data_2 [26]), .Q(n1903) );
  AOI220 U5026 ( .A(n1457), .B(n1409), .C(n1456), .D(n1408), .Q(n4294) );
  NAND21 U5027 ( .A(n4275), .B(n4276), .Q(\execute/old_res [0]) );
  AOI2110 U5028 ( .A(n6512), .B(n6341), .C(n4362), .D(n4363), .Q(n4275) );
  INV0 U5029 ( .A(n3976), .Q(n1442) );
  NOR20 U5030 ( .A(n3692), .B(n4394), .Q(n4134) );
  NOR20 U5031 ( .A(n4394), .B(n3592), .Q(n4270) );
  AOI2110 U5032 ( .A(n1328), .B(n3499), .C(n3679), .D(n3680), .Q(n3678) );
  NOR20 U5033 ( .A(n6341), .B(n4394), .Q(n4400) );
  NOR20 U5034 ( .A(n4394), .B(n5817), .Q(n4355) );
  NAND40 U5035 ( .A(n4176), .B(n4128), .C(n4083), .D(n4111), .Q(n4485) );
  NOR20 U5036 ( .A(n3564), .B(n4394), .Q(n4087) );
  NAND30 U5037 ( .A(n3795), .B(n3757), .C(n3850), .Q(n4513) );
  NOR20 U5038 ( .A(n3542), .B(n6514), .Q(n3543) );
  AOI2110 U5039 ( .A(n6516), .B(n3542), .C(n6512), .D(n3543), .Q(n3541) );
  NAND30 U5040 ( .A(n3436), .B(n3467), .C(n3398), .Q(n4526) );
  AOI210 U5041 ( .A(n6512), .B(n4170), .C(n4102), .Q(n4179) );
  AOI220 U5042 ( .A(n1471), .B(n1422), .C(n6512), .D(n3888), .Q(n3882) );
  AOI2110 U5043 ( .A(n1449), .B(n3886), .C(n1348), .D(n3887), .Q(n3885) );
  AOI220 U5044 ( .A(n1325), .B(n3816), .C(n1321), .D(n3817), .Q(n3809) );
  AOI2110 U5045 ( .A(n6512), .B(n3811), .C(n3812), .D(n3772), .Q(n3810) );
  AOI220 U5046 ( .A(n1325), .B(n3752), .C(n1321), .D(n3838), .Q(n3830) );
  AOI2110 U5047 ( .A(n6512), .B(n3832), .C(n3833), .D(n3772), .Q(n3831) );
  AOI220 U5048 ( .A(n3776), .B(n3777), .C(n1325), .D(n1292), .Q(n3769) );
  AOI220 U5049 ( .A(n1471), .B(n6347), .C(n6512), .D(n3907), .Q(n3902) );
  AOI220 U5050 ( .A(n1347), .B(n3706), .C(n1325), .D(n3496), .Q(n3675) );
  AOI210 U5051 ( .A(n6512), .B(n3757), .C(n3674), .Q(n3748) );
  AOI210 U5052 ( .A(n1321), .B(n3752), .C(n3753), .Q(n3751) );
  AOI220 U5053 ( .A(n3470), .B(n6513), .C(n6512), .D(n3467), .Q(n3458) );
  AOI2110 U5054 ( .A(n1335), .B(n3460), .C(n3461), .D(n3462), .Q(n3459) );
  AOI210 U5055 ( .A(n6512), .B(n3795), .C(n3772), .Q(n3787) );
  AOI210 U5056 ( .A(n1325), .B(n3720), .C(n3791), .Q(n3790) );
  AOI210 U5057 ( .A(n1315), .B(n3713), .C(n3714), .Q(n3712) );
  AOI210 U5058 ( .A(n6512), .B(n3718), .C(n3674), .Q(n3709) );
  AOI220 U5059 ( .A(n3512), .B(n3477), .C(n1331), .D(n3513), .Q(n3489) );
  AOI220 U5060 ( .A(n1328), .B(n3518), .C(n1347), .D(n3519), .Q(n3488) );
  NOR20 U5061 ( .A(n3419), .B(n3398), .Q(n4235) );
  NOR20 U5062 ( .A(n1374), .B(n5830), .Q(n4101) );
  OAI220 U5063 ( .A(n1170), .B(n6063), .C(n1948), .D(n5905), .Q(n2999) );
  OAI220 U5064 ( .A(n1170), .B(n6065), .C(n1948), .D(n5907), .Q(n2936) );
  OAI220 U5065 ( .A(n1170), .B(n6066), .C(n6400), .D(n5840), .Q(n2915) );
  OAI220 U5066 ( .A(n1170), .B(n5939), .C(n1948), .D(n5858), .Q(n2873) );
  OAI220 U5067 ( .A(n1170), .B(n6064), .C(n6401), .D(n5906), .Q(n2957) );
  OAI220 U5068 ( .A(n1162), .B(n6062), .C(n2031), .D(n5904), .Q(n2205) );
  AOI220 U5069 ( .A(n1293), .B(n5830), .C(n1289), .D(n5829), .Q(n4266) );
  AOI220 U5070 ( .A(n6510), .B(n1443), .C(n3616), .D(n6222), .Q(n4267) );
  AOI220 U5071 ( .A(n1293), .B(n6344), .C(n1289), .D(n6345), .Q(n4211) );
  AOI220 U5072 ( .A(n6510), .B(n5830), .C(n3616), .D(n6346), .Q(n4212) );
  AOI220 U5073 ( .A(n1293), .B(n1428), .C(n1289), .D(n6344), .Q(n4268) );
  AOI220 U5074 ( .A(n6510), .B(n6346), .C(n3616), .D(n6345), .Q(n4269) );
  NAND30 U5075 ( .A(n4025), .B(n3998), .C(n3777), .Q(n4500) );
  AOI210 U5076 ( .A(n1446), .B(n3998), .C(n3974), .Q(n3997) );
  OAI310 U5077 ( .A(n6357), .B(n1448), .C(n3907), .D(n3766), .Q(n3906) );
  OAI2110 U5078 ( .A(n3907), .B(n6514), .C(n3918), .D(n3438), .Q(n3904) );
  AOI210 U5079 ( .A(n6512), .B(n3746), .C(n3674), .Q(n3727) );
  AOI220 U5080 ( .A(n1471), .B(n6349), .C(n6512), .D(n3966), .Q(n3959) );
  AOI220 U5081 ( .A(n1470), .B(n1409), .C(n6515), .D(n3746), .Q(n3733) );
  AOI2110 U5082 ( .A(n1335), .B(n3427), .C(n3428), .D(n3429), .Q(n3426) );
  AOI210 U5083 ( .A(n6512), .B(n3436), .C(n3447), .Q(n3424) );
  AOI210 U5084 ( .A(\execute/alu/sll_175/ML_int[4][8] ), .B(n1341), .C(n3444), 
        .Q(n3425) );
  AOI220 U5085 ( .A(\execute/alu/sll_175/ML_int[4][11] ), .B(n1341), .C(n4213), 
        .D(n6513), .Q(n4180) );
  NAND20 U5086 ( .A(n4083), .B(n1439), .Q(n4091) );
  AOI220 U5087 ( .A(n3663), .B(n3657), .C(n1315), .D(n3664), .Q(n3652) );
  AOI220 U5088 ( .A(n6516), .B(n1460), .C(n6515), .D(n3659), .Q(n3666) );
  NAND20 U5089 ( .A(n3662), .B(n3660), .Q(n3665) );
  AOI210 U5090 ( .A(n1305), .B(n3672), .C(n1403), .Q(n3722) );
  OAI2110 U5091 ( .A(n3667), .B(n3744), .C(n3763), .D(n3742), .Q(n3761) );
  NAND20 U5092 ( .A(n1399), .B(n3641), .Q(n3824) );
  AOI220 U5093 ( .A(n3820), .B(n3821), .C(n3822), .D(n6513), .Q(n3807) );
  NOR20 U5094 ( .A(n4083), .B(n3404), .Q(n4084) );
  AOI2110 U5095 ( .A(n3402), .B(n4083), .C(n4084), .D(n6512), .Q(n4081) );
  AOI210 U5096 ( .A(n3851), .B(n3850), .C(n3846), .Q(n3869) );
  AOI220 U5097 ( .A(n3841), .B(n6513), .C(n3842), .D(n3843), .Q(n3828) );
  AOI220 U5098 ( .A(n1293), .B(n6345), .C(n1289), .D(n6346), .Q(n4348) );
  AOI220 U5099 ( .A(n6509), .B(n5829), .C(n6506), .D(n5830), .Q(n4349) );
  AOI220 U5100 ( .A(n1293), .B(n6347), .C(n1289), .D(n1422), .Q(n4396) );
  AOI220 U5101 ( .A(n6509), .B(n1425), .C(n6506), .D(n6193), .Q(n4397) );
  AOI220 U5102 ( .A(n1293), .B(n6346), .C(n1289), .D(n5830), .Q(n4144) );
  AOI220 U5103 ( .A(n3615), .B(n6222), .C(n6507), .D(n5829), .Q(n4145) );
  AOI220 U5104 ( .A(n1293), .B(n5829), .C(n1289), .D(n6222), .Q(n4207) );
  AOI220 U5105 ( .A(n6510), .B(n1445), .C(n6506), .D(n1443), .Q(n4208) );
  NOR20 U5106 ( .A(n4170), .B(n6514), .Q(n4197) );
  AOI2110 U5107 ( .A(n6516), .B(n4170), .C(n4197), .D(n6512), .Q(n4196) );
  AOI220 U5108 ( .A(n1293), .B(n1426), .C(n1289), .D(n1427), .Q(n4346) );
  AOI220 U5109 ( .A(n6509), .B(n6344), .C(n6506), .D(n1428), .Q(n4347) );
  OAI2110 U5110 ( .A(n3467), .B(n6514), .C(n3468), .D(n6352), .Q(n3466) );
  AOI220 U5111 ( .A(n3464), .B(n3465), .C(n3466), .D(n1425), .Q(n3463) );
  NAND20 U5112 ( .A(n3742), .B(n3741), .Q(n3785) );
  NOR20 U5113 ( .A(n1454), .B(n3777), .Q(n3783) );
  AOI220 U5114 ( .A(n1470), .B(n1367), .C(n6515), .D(n4170), .Q(n4200) );
  OAI310 U5115 ( .A(n3407), .B(n1298), .C(n4165), .D(n3438), .Q(n4163) );
  AOI210 U5116 ( .A(n3599), .B(n3600), .C(n3601), .Q(n3598) );
  AOI220 U5117 ( .A(n1293), .B(n1427), .C(n1289), .D(n1428), .Q(n3955) );
  OAI310 U5118 ( .A(n4225), .B(n4226), .C(n6512), .D(n4176), .Q(n4224) );
  NOR20 U5119 ( .A(n3998), .B(n3404), .Q(n4007) );
  AOI2110 U5120 ( .A(n3402), .B(n3998), .C(n4007), .D(n6512), .Q(n4004) );
  AOI220 U5121 ( .A(n3878), .B(n1218), .C(\execute/alu/sll_175/ML_int[3][18] ), 
        .D(n3507), .Q(n4005) );
  NOR20 U5122 ( .A(n3850), .B(n3404), .Q(n3879) );
  AOI2110 U5123 ( .A(n3402), .B(n3850), .C(n3879), .D(n6512), .Q(n3876) );
  AOI220 U5124 ( .A(n3878), .B(\execute/alu/sll_175/ML_int[3][6] ), .C(
        \execute/alu/sll_175/ML_int[3][22] ), .D(n3507), .Q(n3877) );
  NAND20 U5125 ( .A(n3662), .B(n3657), .Q(n3635) );
  AOI310 U5126 ( .A(n1341), .B(n5819), .C(\execute/alu/sll_175/ML_int[3][10] ), 
        .D(n1348), .Q(n4009) );
  AOI220 U5127 ( .A(n1470), .B(n1385), .C(n6515), .D(n3998), .Q(n4008) );
  OAI310 U5128 ( .A(n3407), .B(n4129), .C(n4130), .D(n3438), .Q(n4126) );
  INV0 U5129 ( .A(n3477), .Q(n1358) );
  INV0 U5130 ( .A(n3436), .Q(n1361) );
  INV0 U5131 ( .A(n3657), .Q(n1411) );
  AOI220 U5132 ( .A(n6356), .B(n5829), .C(n1258), .D(n6346), .Q(n4143) );
  AOI220 U5133 ( .A(n1372), .B(n6346), .C(n1374), .D(n5830), .Q(n4315) );
  OAI220 U5134 ( .A(n3998), .B(n3999), .C(n4025), .D(n4018), .Q(n4339) );
  AOI220 U5135 ( .A(n4025), .B(n4018), .C(n4024), .D(n4039), .Q(n4340) );
  AOI220 U5136 ( .A(n3602), .B(n6345), .C(n1258), .D(n1428), .Q(n4258) );
  OAI310 U5137 ( .A(n6357), .B(n5829), .C(n4083), .D(n3766), .Q(n4072) );
  NOR20 U5138 ( .A(n6341), .B(n1310), .Q(n3602) );
  NOR20 U5139 ( .A(n3476), .B(n3477), .Q(n3473) );
  OAI210 U5140 ( .A(n3473), .B(n3474), .C(n6250), .Q(n3472) );
  AOI220 U5141 ( .A(n1470), .B(n1387), .C(n6515), .D(n3966), .Q(n3965) );
  CLKIN1 U5142 ( .A(n6960), .Q(n6959) );
  CLKIN1 U5143 ( .A(n6984), .Q(n6983) );
  CLKIN1 U5144 ( .A(n6978), .Q(n6977) );
  CLKIN1 U5145 ( .A(n6952), .Q(n6951) );
  CLKIN1 U5146 ( .A(n6994), .Q(n6993) );
  CLKIN1 U5147 ( .A(n6974), .Q(n6973) );
  CLKIN1 U5148 ( .A(n6972), .Q(n6971) );
  CLKIN1 U5149 ( .A(n6970), .Q(n6969) );
  CLKIN1 U5150 ( .A(n6966), .Q(n6965) );
  CLKIN1 U5151 ( .A(n6956), .Q(n6955) );
  CLKIN1 U5152 ( .A(n6938), .Q(n6937) );
  NAND20 U5153 ( .A(n1310), .B(n6341), .Q(n4131) );
  BUF2 U5154 ( .A(inst_out[25]), .Q(n6498) );
  BUF2 U5155 ( .A(inst_out[20]), .Q(n6492) );
  AOI220 U5156 ( .A(n1415), .B(n1258), .C(n6349), .D(n6356), .Q(n3944) );
  AOI210 U5157 ( .A(n3944), .B(n3945), .C(n3601), .Q(n3943) );
  OAI2110 U5158 ( .A(n6349), .B(n3583), .C(n3504), .D(n3584), .Q(n3581) );
  AOI220 U5159 ( .A(n3585), .B(n6349), .C(n3586), .D(n6513), .Q(n3584) );
  NAND30 U5160 ( .A(n6321), .B(n4343), .C(n4064), .Q(n3399) );
  AOI220 U5161 ( .A(n1258), .B(n5829), .C(n6355), .D(n1445), .Q(n4190) );
  AOI220 U5162 ( .A(n6356), .B(n1422), .C(n1258), .D(n6349), .Q(n3600) );
  AOI220 U5163 ( .A(n6355), .B(n6349), .C(n1294), .D(n1415), .Q(n4370) );
  AOI210 U5164 ( .A(n4370), .B(n4371), .C(n3601), .Q(n4369) );
  OAI220 U5165 ( .A(n3811), .B(n3821), .C(n3832), .D(n3843), .Q(n4300) );
  AOI220 U5166 ( .A(n3832), .B(n3843), .C(n3850), .D(n3870), .Q(n4299) );
  AOI220 U5167 ( .A(n3811), .B(n3821), .C(n3795), .D(n3793), .Q(n4302) );
  AOI220 U5168 ( .A(n6355), .B(n1422), .C(n1294), .D(n6349), .Q(n3701) );
  NOR20 U5169 ( .A(n6204), .B(n3692), .Q(n3689) );
  AOI220 U5170 ( .A(n6355), .B(n5830), .C(n1258), .D(n6344), .Q(n4205) );
  AOI220 U5171 ( .A(n3602), .B(n5830), .C(n1258), .D(n6345), .Q(n4374) );
  AOI220 U5172 ( .A(n6356), .B(n1428), .C(n1258), .D(n1426), .Q(n4379) );
  AOI220 U5173 ( .A(n6356), .B(n6344), .C(n1258), .D(n1427), .Q(n3947) );
  NAND20 U5174 ( .A(n3936), .B(n3937), .Q(n3693) );
  AOI220 U5175 ( .A(n3602), .B(n6222), .C(n1258), .D(n5830), .Q(n4253) );
  AOI220 U5176 ( .A(n6355), .B(n1425), .C(n1294), .D(n1422), .Q(n4376) );
  AOI220 U5177 ( .A(n6356), .B(n6193), .C(n1258), .D(n6347), .Q(n4377) );
  NOR20 U5178 ( .A(n4282), .B(n1476), .Q(n4064) );
  NAND20 U5179 ( .A(n1320), .B(n3592), .Q(n3605) );
  NOR20 U5180 ( .A(n5946), .B(n1992), .Q(n1989) );
  OAI2110 U5181 ( .A(n3888), .B(n6514), .C(n3889), .D(n3438), .Q(n3886) );
  NAND20 U5182 ( .A(n6516), .B(n3888), .Q(n3889) );
  OAI2110 U5183 ( .A(n3436), .B(n6514), .C(n3437), .D(n6352), .Q(n3435) );
  NAND20 U5184 ( .A(n6516), .B(n3436), .Q(n3437) );
  NOR30 U5185 ( .A(n4395), .B(n6321), .C(n4343), .Q(n4068) );
  AOI220 U5186 ( .A(n1470), .B(n1396), .C(n6515), .D(n3850), .Q(n3880) );
  AOI2110 U5187 ( .A(n3402), .B(n4111), .C(n4112), .D(n6512), .Q(n4107) );
  NOR20 U5188 ( .A(n4111), .B(n3404), .Q(n4112) );
  OAI220 U5189 ( .A(n1356), .B(n6514), .C(n3542), .D(n6358), .Q(n3537) );
  OAI220 U5190 ( .A(n1360), .B(n3404), .C(n3467), .D(n6358), .Q(n3464) );
  NOR20 U5191 ( .A(n3718), .B(n3404), .Q(n3719) );
  AOI2110 U5192 ( .A(n3402), .B(n3718), .C(n3719), .D(n6512), .Q(n3715) );
  AOI220 U5193 ( .A(n1470), .B(n1410), .C(n6515), .D(n3718), .Q(n3717) );
  NOR20 U5194 ( .A(n3795), .B(n6514), .Q(n3796) );
  AOI2110 U5195 ( .A(n3402), .B(n3795), .C(n3796), .D(n6512), .Q(n3792) );
  AOI220 U5196 ( .A(n1470), .B(n1404), .C(n6515), .D(n3795), .Q(n3794) );
  NOR20 U5197 ( .A(n3757), .B(n3404), .Q(n3758) );
  AOI2110 U5198 ( .A(n3402), .B(n3757), .C(n3758), .D(n6512), .Q(n3754) );
  AOI220 U5199 ( .A(n1470), .B(n1408), .C(n6515), .D(n3757), .Q(n3756) );
  NAND20 U5200 ( .A(n1338), .B(n5817), .Q(n4372) );
  AOI210 U5201 ( .A(n6515), .B(n1259), .C(n4344), .Q(n4341) );
  AOI220 U5202 ( .A(n1470), .B(n1259), .C(n6515), .D(n6341), .Q(n4342) );
  XNR20 U5203 ( .A(n6351), .B(n4380), .Q(n4364) );
  OAI2110 U5204 ( .A(n3811), .B(n6514), .C(n3819), .D(n6352), .Q(n3818) );
  NAND20 U5205 ( .A(n6516), .B(n3811), .Q(n3819) );
  OAI2110 U5206 ( .A(n3832), .B(n6514), .C(n3840), .D(n6352), .Q(n3839) );
  NAND20 U5207 ( .A(n6516), .B(n3832), .Q(n3840) );
  OAI2110 U5208 ( .A(n3746), .B(n6514), .C(n3747), .D(n3438), .Q(n3730) );
  NAND20 U5209 ( .A(n6516), .B(n3746), .Q(n3747) );
  OAI2110 U5210 ( .A(n3966), .B(n6514), .C(n3978), .D(n6352), .Q(n3962) );
  NAND20 U5211 ( .A(n3402), .B(n3966), .Q(n3978) );
  NOR20 U5212 ( .A(n3777), .B(n3404), .Q(n3782) );
  NOR30 U5213 ( .A(n6357), .B(n1449), .C(n3888), .Q(n3887) );
  NOR30 U5214 ( .A(n6357), .B(n1460), .C(n3657), .Q(n3656) );
  OAI220 U5215 ( .A(n1310), .B(n3404), .C(n3692), .D(n6358), .Q(n3949) );
  OAI210 U5216 ( .A(n4025), .B(n6514), .C(n6352), .Q(n4013) );
  INV0 U5217 ( .A(n6349), .Q(n1418) );
  INV0 U5218 ( .A(n3850), .Q(n1396) );
  NAND20 U5219 ( .A(n6516), .B(n3467), .Q(n3468) );
  NAND20 U5220 ( .A(n6516), .B(n3907), .Q(n3918) );
  INV0 U5221 ( .A(\execute/op_21 [30]), .Q(n1459) );
  INV0 U5222 ( .A(n3564), .Q(n1344) );
  NOR30 U5223 ( .A(n6351), .B(n4395), .C(n4343), .Q(n4366) );
  XNR20 U5224 ( .A(write_register[4]), .B(rs[4]), .Q(n4546) );
  NAND42 U5225 ( .A(n4545), .B(n4546), .C(n4547), .D(n4548), .Q(n4542) );
  XNR20 U5226 ( .A(write_register[3]), .B(rs[3]), .Q(n4547) );
  XNR20 U5227 ( .A(rs[1]), .B(n5848), .Q(n4551) );
  XNR20 U5228 ( .A(rs[2]), .B(n5941), .Q(n4550) );
  NOR30 U5229 ( .A(n1494), .B(n1461), .C(n1991), .Q(n1990) );
  AOI220 U5230 ( .A(ram_adr[24]), .B(n6337), .C(n6339), .D(data_1[24]), .Q(
        n4517) );
  AOI220 U5231 ( .A(n6503), .B(n6979), .C(pc_ex[24]), .D(n6323), .Q(n4516) );
  AOI220 U5232 ( .A(n6503), .B(n6943), .C(pc_ex[6]), .D(n6324), .Q(n4518) );
  AOI220 U5233 ( .A(ram_adr[6]), .B(n6336), .C(n6339), .D(data_1[6]), .Q(n4519) );
  AOI220 U5234 ( .A(n6503), .B(write_data_reg[27]), .C(pc_ex[27]), .D(n6324), 
        .Q(n4522) );
  AOI220 U5235 ( .A(ram_adr[25]), .B(n6337), .C(n6339), .D(data_1[25]), .Q(
        n4525) );
  AOI220 U5236 ( .A(n6503), .B(write_data_reg[25]), .C(pc_ex[25]), .D(n6323), 
        .Q(n4524) );
  AOI220 U5237 ( .A(ram_adr[14]), .B(n6336), .C(n6340), .D(data_1[14]), .Q(
        n4493) );
  AOI220 U5238 ( .A(n6503), .B(write_data_reg[30]), .C(pc_ex[30]), .D(n6324), 
        .Q(n4527) );
  AOI220 U5239 ( .A(ram_adr[26]), .B(n6337), .C(n6340), .D(data_1[26]), .Q(
        n4508) );
  AOI220 U5240 ( .A(ram_adr[21]), .B(n6337), .C(n6340), .D(data_1[21]), .Q(
        n4504) );
  AOI220 U5241 ( .A(n6503), .B(write_data_reg[21]), .C(pc_ex[21]), .D(n6323), 
        .Q(n4503) );
  AOI220 U5242 ( .A(ram_adr[28]), .B(n6337), .C(n6339), .D(data_1[28]), .Q(
        n4530) );
  AOI220 U5243 ( .A(n6503), .B(write_data_reg[28]), .C(pc_ex[28]), .D(n6324), 
        .Q(n4529) );
  AOI220 U5244 ( .A(ram_adr[17]), .B(n6337), .C(n6339), .D(data_1[17]), .Q(
        n4512) );
  AOI220 U5245 ( .A(n6503), .B(write_data_reg[17]), .C(pc_ex[17]), .D(n6323), 
        .Q(n4511) );
  AOI220 U5246 ( .A(ram_adr[16]), .B(n6336), .C(n6340), .D(data_1[16]), .Q(
        n4506) );
  AOI220 U5247 ( .A(n6503), .B(n6963), .C(pc_ex[16]), .D(n6324), .Q(n4505) );
  AOI220 U5248 ( .A(n6504), .B(write_data_reg[10]), .C(pc_ex[10]), .D(n6323), 
        .Q(n4498) );
  AOI220 U5249 ( .A(ram_adr[10]), .B(n6337), .C(n6340), .D(data_1[10]), .Q(
        n4499) );
  AOI220 U5250 ( .A(n6504), .B(n6957), .C(pc_ex[13]), .D(n6324), .Q(n4496) );
  AOI220 U5251 ( .A(ram_adr[13]), .B(n6336), .C(n6340), .D(data_1[13]), .Q(
        n4497) );
  AOI220 U5252 ( .A(n1827), .B(n6314), .C(n1142), .D(inst_out[23]), .Q(n1826)
         );
  NOR20 U5253 ( .A(n6286), .B(n1137), .Q(n5763) );
  NOR20 U5254 ( .A(n6286), .B(n1117), .Q(n5743) );
  AOI220 U5255 ( .A(n1792), .B(n6314), .C(n1142), .D(inst_out[21]), .Q(n1791)
         );
  AOI220 U5256 ( .A(n1786), .B(n6315), .C(n1142), .D(inst_out[17]), .Q(n1785)
         );
  CLKIN3 U5257 ( .A(\execute/op_21 [15]), .Q(n1440) );
  AOI220 U5258 ( .A(n6504), .B(n6941), .C(pc_ex[5]), .D(n6323), .Q(n4402) );
  AOI220 U5259 ( .A(ram_adr[5]), .B(n6337), .C(n6340), .D(data_1[5]), .Q(n4403) );
  OAI310 U5260 ( .A(n5946), .B(n5627), .C(n4409), .D(n4410), .Q(n4407) );
  AOI220 U5261 ( .A(n6504), .B(write_data_reg[12]), .C(pc_ex[12]), .D(n6324), 
        .Q(n4488) );
  AOI220 U5262 ( .A(ram_adr[12]), .B(n6336), .C(n6340), .D(data_1[12]), .Q(
        n4489) );
  AOI220 U5263 ( .A(ram_adr[31]), .B(n6336), .C(n6339), .D(data_1[31]), .Q(
        n4540) );
  AOI220 U5264 ( .A(n6503), .B(write_data_reg[31]), .C(pc_ex[31]), .D(n6324), 
        .Q(n4539) );
  AOI220 U5265 ( .A(n6332), .B(data_2[12]), .C(n5815), .D(ram_adr[12]), .Q(
        n4455) );
  AOI220 U5266 ( .A(n6333), .B(data_2[22]), .C(n5816), .D(ram_adr[22]), .Q(
        n4443) );
  AOI220 U5267 ( .A(n6332), .B(data_2[20]), .C(n5816), .D(ram_adr[20]), .Q(
        n4446) );
  AOI220 U5268 ( .A(n1467), .B(n6074), .C(pc_ex[2]), .D(n6324), .Q(n4466) );
  AOI220 U5269 ( .A(n6330), .B(data_2[8]), .C(n5816), .D(ram_adr[8]), .Q(n4429) );
  AOI220 U5270 ( .A(n6332), .B(data_2[15]), .C(n5816), .D(ram_adr[15]), .Q(
        n4452) );
  AOI220 U5271 ( .A(n6333), .B(data_2[21]), .C(n5816), .D(ram_adr[21]), .Q(
        n4445) );
  AOI220 U5272 ( .A(n6330), .B(data_2[27]), .C(n5816), .D(ram_adr[27]), .Q(
        n4438) );
  CLKIN6 U5273 ( .A(rt[3]), .Q(n1489) );
  XNR20 U5274 ( .A(write_register[2]), .B(rt[2]), .Q(n4561) );
  INV2 U5275 ( .A(n1971), .Q(n1150) );
  NAND30 U5276 ( .A(n6279), .B(n1972), .C(n5716), .Q(n1971) );
  INV0 U5277 ( .A(\wb_WB[0] ), .Q(n6929) );
  AOI220 U5278 ( .A(ram_adr[4]), .B(n6336), .C(n6340), .D(data_1[4]), .Q(n4459) );
  AOI220 U5279 ( .A(n1467), .B(n6073), .C(pc_ex[4]), .D(n6324), .Q(n4460) );
  AOI220 U5280 ( .A(n6364), .B(n5940), .C(n6370), .D(n5426), .Q(n3168) );
  OAI221 U5281 ( .A(n4691), .B(n6415), .C(n4690), .D(n6417), .Q(n1916) );
  OAI221 U5282 ( .A(n4679), .B(n6479), .C(n4678), .D(n6481), .Q(n2526) );
  OAI221 U5283 ( .A(n4663), .B(n6415), .C(n4662), .D(n6417), .Q(n3131) );
  OAI221 U5284 ( .A(n4623), .B(n6479), .C(n4622), .D(n6481), .Q(n2400) );
  OAI221 U5285 ( .A(n4703), .B(n6479), .C(n4702), .D(n6481), .Q(n2652) );
  OAI221 U5286 ( .A(n4667), .B(n6479), .C(n4666), .D(n6481), .Q(n2463) );
  OAI221 U5287 ( .A(n4615), .B(n6478), .C(n4614), .D(n6480), .Q(n2358) );
  OAI221 U5288 ( .A(n4695), .B(n6478), .C(n4694), .D(n6480), .Q(n2610) );
  OAI221 U5289 ( .A(n4683), .B(n6478), .C(n4682), .D(n6480), .Q(n2547) );
  OAI221 U5290 ( .A(n4603), .B(n6478), .C(n4602), .D(n6480), .Q(n2295) );
  OAI221 U5291 ( .A(n4627), .B(n6478), .C(n4626), .D(n6480), .Q(n2421) );
  OAI221 U5292 ( .A(n4587), .B(n2022), .C(n4586), .D(n2023), .Q(n2190) );
  OAI221 U5293 ( .A(n4671), .B(n1939), .C(n4670), .D(n1940), .Q(n3173) );
  OAI221 U5294 ( .A(n4675), .B(n2022), .C(n4674), .D(n2023), .Q(n2505) );
  OAI221 U5295 ( .A(n4687), .B(n2022), .C(n4686), .D(n2023), .Q(n2568) );
  OAI221 U5296 ( .A(n4619), .B(n2022), .C(n4618), .D(n2023), .Q(n2379) );
  OAI221 U5297 ( .A(n4699), .B(n2022), .C(n4698), .D(n2023), .Q(n2631) );
  OAI221 U5298 ( .A(n4639), .B(n2022), .C(n4638), .D(n2023), .Q(n2064) );
  AOI220 U5299 ( .A(n6332), .B(data_2[30]), .C(n5816), .D(ram_adr[30]), .Q(
        n4434) );
  AOI220 U5300 ( .A(n1467), .B(n6075), .C(pc_ex[3]), .D(n6323), .Q(n4462) );
  NOR42 U5301 ( .A(n2989), .B(n2990), .C(n2991), .D(n2992), .Q(n2988) );
  NOR41 U5302 ( .A(n2993), .B(n2994), .C(n2995), .D(n2996), .Q(n2987) );
  NOR41 U5303 ( .A(n2947), .B(n2948), .C(n2949), .D(n2950), .Q(n2946) );
  AOI220 U5304 ( .A(n6329), .B(data_2[18]), .C(n5815), .D(ram_adr[18]), .Q(
        n4449) );
  AOI220 U5305 ( .A(n6329), .B(data_2[28]), .C(n5816), .D(ram_adr[28]), .Q(
        n4437) );
  AOI220 U5306 ( .A(n6333), .B(data_2[24]), .C(n5815), .D(ram_adr[24]), .Q(
        n4441) );
  AOI220 U5307 ( .A(n6332), .B(data_2[29]), .C(n5815), .D(ram_adr[29]), .Q(
        n4436) );
  AOI220 U5308 ( .A(n6330), .B(data_2[25]), .C(n5816), .D(ram_adr[25]), .Q(
        n4440) );
  AOI220 U5309 ( .A(n6329), .B(data_2[26]), .C(n5815), .D(ram_adr[26]), .Q(
        n4439) );
  AOI220 U5310 ( .A(n6330), .B(data_2[19]), .C(n5816), .D(ram_adr[19]), .Q(
        n4448) );
  AOI310 U5311 ( .A(n5696), .B(n4414), .C(n1493), .D(n6233), .Q(n4411) );
  OAI2110 U5312 ( .A(n4411), .B(n5999), .C(n1481), .D(n4412), .Q(n4282) );
  CLKIN1 U5313 ( .A(n5734), .Q(n6490) );
  NAND20 U5314 ( .A(n4409), .B(n5627), .Q(n4420) );
  OAI310 U5315 ( .A(n4415), .B(n6216), .C(n4408), .D(n4416), .Q(n4281) );
  OAI2110 U5316 ( .A(n6246), .B(n5946), .C(n4420), .D(n5696), .Q(n4415) );
  OAI210 U5317 ( .A(n5694), .B(n5999), .C(n1986), .Q(n4343) );
  AOI220 U5318 ( .A(n6330), .B(data_2[31]), .C(n5815), .D(ram_adr[31]), .Q(
        n4559) );
  NAND30 U5319 ( .A(n5867), .B(n5941), .C(write_register[1]), .Q(n1958) );
  NAND30 U5320 ( .A(write_register[2]), .B(n5867), .C(write_register[1]), .Q(
        n1962) );
  NAND30 U5321 ( .A(n5867), .B(n5848), .C(write_register[2]), .Q(n1956) );
  XNR20 U5322 ( .A(rt[2]), .B(n5727), .Q(n3384) );
  XNR20 U5323 ( .A(rt[2]), .B(n5726), .Q(n3378) );
  XNR20 U5324 ( .A(n1485), .B(n5728), .Q(n3380) );
  XNR20 U5325 ( .A(n6209), .B(n5724), .Q(n3381) );
  XNR20 U5326 ( .A(n1485), .B(n5725), .Q(n3386) );
  XNR20 U5327 ( .A(n6209), .B(n5723), .Q(n3387) );
  AOI220 U5328 ( .A(data_1[30]), .B(n6339), .C(n6336), .D(ram_adr[30]), .Q(
        n4289) );
  OAI220 U5329 ( .A(n4364), .B(n3407), .C(n4365), .D(n3596), .Q(n4363) );
  INV3 U5330 ( .A(n6352), .Q(n6512) );
  INV3 U5331 ( .A(n6312), .Q(n6288) );
  INV3 U5332 ( .A(n6312), .Q(n6281) );
  INV3 U5333 ( .A(n3570), .Q(n1321) );
  INV3 U5334 ( .A(n3554), .Q(n1328) );
  NOR21 U5335 ( .A(n3948), .B(n5819), .Q(n5811) );
  INV3 U5336 ( .A(n3534), .Q(n1325) );
  INV3 U5337 ( .A(n3540), .Q(n1331) );
  BUF2 U5338 ( .A(n3438), .Q(n6352) );
  INV3 U5339 ( .A(n3667), .Q(n1306) );
  INV3 U5340 ( .A(n3743), .Q(n1305) );
  AOI221 U5341 ( .A(n1341), .B(n5809), .C(n3530), .D(n1321), .Q(n3529) );
  AOI221 U5342 ( .A(n3647), .B(n1342), .C(n6343), .D(n6258), .Q(n3644) );
  NAND22 U5343 ( .A(n3649), .B(n6756), .Q(n3648) );
  NAND22 U5344 ( .A(\execute/alu/sll_175/ML_int[3][4] ), .B(n6756), .Q(n1856)
         );
  NOR21 U5345 ( .A(n1222), .B(n5819), .Q(n5809) );
  INV3 U5346 ( .A(\execute/alu/sll_175/ML_int[3][5] ), .Q(n1222) );
  INV3 U5347 ( .A(n4129), .Q(n1299) );
  INV3 U5348 ( .A(n4464), .Q(n1218) );
  NAND22 U5349 ( .A(\execute/alu/sll_175/ML_int[2][2] ), .B(n6759), .Q(n4464)
         );
  INV3 U5350 ( .A(n3778), .Q(n1304) );
  NAND22 U5351 ( .A(\execute/alu/sll_175/ML_int[3][7] ), .B(n6756), .Q(n3487)
         );
  IMUX21 U5352 ( .A(\execute/alu/sll_175/ML_int[3][20] ), .B(
        \execute/alu/sll_175/ML_int[3][12] ), .S(n5819), .Q(n6259) );
  NAND22 U5353 ( .A(n1473), .B(n3454), .Q(n3570) );
  NAND22 U5354 ( .A(n1473), .B(n3455), .Q(n3534) );
  NAND22 U5355 ( .A(n1473), .B(n1329), .Q(n3554) );
  INV3 U5356 ( .A(n6759), .Q(n6758) );
  INV3 U5357 ( .A(n4262), .Q(n1273) );
  NAND22 U5358 ( .A(n1473), .B(n1332), .Q(n3540) );
  INV3 U5359 ( .A(n3430), .Q(n1333) );
  INV3 U5360 ( .A(n3535), .Q(n1335) );
  INV3 U5361 ( .A(n3431), .Q(n1313) );
  NAND22 U5362 ( .A(n1224), .B(n6756), .Q(n1855) );
  AOI221 U5363 ( .A(n3859), .B(n3706), .C(n6236), .D(n3705), .Q(n3989) );
  INV3 U5364 ( .A(n3995), .Q(n1292) );
  INV3 U5365 ( .A(n3414), .Q(n1332) );
  NOR21 U5366 ( .A(n1226), .B(n5820), .Q(n5810) );
  INV3 U5367 ( .A(\execute/alu/sll_175/ML_int[1][1] ), .Q(n1226) );
  NOR21 U5368 ( .A(n1214), .B(n6757), .Q(n5808) );
  INV3 U5369 ( .A(n3838), .Q(n1280) );
  INV3 U5370 ( .A(n6343), .Q(n1342) );
  INV3 U5371 ( .A(n3415), .Q(n1329) );
  INV3 U5372 ( .A(n6511), .Q(n6509) );
  INV3 U5373 ( .A(n3817), .Q(n1266) );
  INV3 U5374 ( .A(n3797), .Q(n1286) );
  INV3 U5375 ( .A(n3455), .Q(n1326) );
  INV3 U5376 ( .A(n3557), .Q(n1263) );
  INV3 U5377 ( .A(n3544), .Q(n1283) );
  IMUX21 U5378 ( .A(\execute/alu/sll_175/ML_int[3][19] ), .B(
        \execute/alu/sll_175/ML_int[3][11] ), .S(n5819), .Q(n6260) );
  NAND22 U5379 ( .A(n1347), .B(n1323), .Q(n4105) );
  INV3 U5380 ( .A(n3553), .Q(n1347) );
  INV3 U5381 ( .A(n3859), .Q(n1346) );
  INV3 U5382 ( .A(n3453), .Q(n1339) );
  INV3 U5383 ( .A(n3982), .Q(n1245) );
  INV3 U5384 ( .A(n6517), .Q(n6516) );
  INV3 U5385 ( .A(n6373), .Q(n6375) );
  INV3 U5386 ( .A(n6373), .Q(n6374) );
  INV3 U5387 ( .A(n6435), .Q(n6436) );
  INV3 U5388 ( .A(n6373), .Q(n6376) );
  INV3 U5389 ( .A(n6435), .Q(n6437) );
  INV3 U5390 ( .A(n6435), .Q(n6438) );
  INV3 U5391 ( .A(n3504), .Q(n1354) );
  INV3 U5392 ( .A(n3814), .Q(n1227) );
  INV3 U5393 ( .A(n3759), .Q(n1240) );
  INV3 U5394 ( .A(n3575), .Q(n1231) );
  INV3 U5395 ( .A(n6373), .Q(n6377) );
  INV3 U5396 ( .A(n6435), .Q(n6439) );
  AOI211 U5397 ( .A(n3802), .B(n6213), .C(n3803), .Q(n3667) );
  BUF2 U5398 ( .A(n1777), .Q(n6487) );
  BUF2 U5399 ( .A(n1777), .Q(n6488) );
  INV3 U5400 ( .A(n3601), .Q(n1317) );
  NAND22 U5401 ( .A(n3914), .B(n3912), .Q(n3637) );
  INV3 U5402 ( .A(n6505), .Q(n6504) );
  INV3 U5403 ( .A(n3899), .Q(n1390) );
  INV3 U5404 ( .A(n3591), .Q(n1319) );
  INV3 U5405 ( .A(n1868), .Q(n1160) );
  NAND41 U5406 ( .A(n4154), .B(n4155), .C(n4156), .D(n4157), .Q(
        \execute/old_res [12]) );
  NAND41 U5407 ( .A(n4113), .B(n4114), .C(n4115), .D(n4116), .Q(
        \execute/old_res [13]) );
  NAND41 U5408 ( .A(n4093), .B(n4094), .C(n4095), .D(n4096), .Q(
        \execute/old_res [14]) );
  NOR31 U5409 ( .A(n4097), .B(n4098), .C(n4099), .Q(n4096) );
  AOI211 U5410 ( .A(n1471), .B(n1427), .C(n3798), .Q(n3788) );
  NAND22 U5411 ( .A(n1402), .B(n3764), .Q(n3801) );
  NAND22 U5412 ( .A(n1461), .B(n1258), .Q(n3624) );
  AOI221 U5413 ( .A(n1321), .B(n3775), .C(\execute/alu/sll_175/ML_int[5][26] ), 
        .D(n1353), .Q(n3774) );
  NAND22 U5414 ( .A(n3741), .B(n3764), .Q(n3744) );
  INV3 U5415 ( .A(n4003), .Q(n1382) );
  NAND22 U5416 ( .A(n3871), .B(n1391), .Q(n3897) );
  AOI211 U5417 ( .A(n3893), .B(n6513), .C(n1248), .Q(n3883) );
  INV3 U5418 ( .A(n3894), .Q(n1248) );
  XNR21 U5419 ( .A(n3897), .B(n3898), .Q(n3893) );
  AOI221 U5420 ( .A(n6515), .B(n3895), .C(n3533), .D(n6236), .Q(n3894) );
  NAND22 U5421 ( .A(n1314), .B(n6236), .Q(n3431) );
  NAND22 U5422 ( .A(n1336), .B(n6236), .Q(n3535) );
  NAND22 U5423 ( .A(n4263), .B(n4264), .Q(n3775) );
  AOI221 U5424 ( .A(n1293), .B(n1454), .C(n1289), .D(n1456), .Q(n4263) );
  AOI221 U5425 ( .A(n6510), .B(n1458), .C(n6506), .D(n1457), .Q(n4264) );
  NAND22 U5426 ( .A(n1334), .B(n6236), .Q(n3430) );
  NAND22 U5427 ( .A(n4273), .B(n4274), .Q(n3867) );
  NAND22 U5428 ( .A(n4201), .B(n4202), .Q(n3752) );
  NOR21 U5429 ( .A(n4069), .B(n3863), .Q(n3454) );
  NOR21 U5430 ( .A(n4069), .B(n3890), .Q(n3455) );
  NAND22 U5431 ( .A(n1473), .B(n4265), .Q(n3553) );
  NAND22 U5432 ( .A(n1327), .B(n4265), .Q(n3417) );
  NAND22 U5433 ( .A(n4353), .B(n4354), .Q(n3816) );
  NAND22 U5434 ( .A(n4360), .B(n4361), .Q(n3557) );
  NAND22 U5435 ( .A(n4356), .B(n4357), .Q(n3817) );
  NAND22 U5436 ( .A(n1323), .B(n4265), .Q(n3416) );
  AOI221 U5437 ( .A(n3532), .B(n1315), .C(n3533), .D(n1349), .Q(n3531) );
  AOI221 U5438 ( .A(n3981), .B(n1335), .C(n3837), .D(n1333), .Q(n4092) );
  NAND22 U5439 ( .A(n4150), .B(n4151), .Q(n3544) );
  NAND22 U5440 ( .A(n4121), .B(n4122), .Q(n3797) );
  AOI221 U5441 ( .A(n6509), .B(n1457), .C(n6507), .D(n1456), .Q(n4122) );
  OAI2111 U5442 ( .A(n1286), .B(n3890), .C(n3864), .D(n3891), .Q(n3546) );
  NAND22 U5443 ( .A(n3994), .B(n1345), .Q(n3414) );
  INV3 U5444 ( .A(n3569), .Q(n1341) );
  OAI2111 U5445 ( .A(n1270), .B(n3863), .C(n3864), .D(n3865), .Q(n3519) );
  AOI221 U5446 ( .A(n1292), .B(n3866), .C(n1327), .D(n3775), .Q(n3865) );
  NAND22 U5447 ( .A(n3866), .B(n1345), .Q(n3415) );
  OAI2111 U5448 ( .A(n1280), .B(n3890), .C(n3864), .D(n3977), .Q(n3580) );
  AOI221 U5449 ( .A(n1323), .B(n3485), .C(n3866), .D(n3752), .Q(n3977) );
  BUF2 U5450 ( .A(\execute/alu/sll_175/temp_int_SH[4] ), .Q(n6343) );
  NAND22 U5451 ( .A(n4351), .B(n4352), .Q(n4066) );
  NAND22 U5452 ( .A(n4198), .B(n4199), .Q(n3838) );
  NOR21 U5453 ( .A(n4350), .B(n1359), .Q(n4067) );
  NAND22 U5454 ( .A(n3992), .B(n3993), .Q(n3706) );
  AOI221 U5455 ( .A(n1327), .B(n3867), .C(n1323), .D(n3513), .Q(n3993) );
  NAND22 U5456 ( .A(n3613), .B(n3614), .Q(n3482) );
  NAND22 U5457 ( .A(n3707), .B(n3708), .Q(n3496) );
  NOR21 U5458 ( .A(n1216), .B(n5820), .Q(\execute/alu/sll_175/ML_int[2][0] )
         );
  INV3 U5459 ( .A(n3890), .Q(n1327) );
  NAND22 U5460 ( .A(n3957), .B(n3958), .Q(n3530) );
  NAND22 U5461 ( .A(n4026), .B(n4027), .Q(n3954) );
  INV3 U5462 ( .A(n3615), .Q(n6511) );
  INV3 U5463 ( .A(n3616), .Q(n6508) );
  INV3 U5464 ( .A(n3720), .Q(n1288) );
  INV3 U5465 ( .A(n4069), .Q(n1345) );
  INV3 U5466 ( .A(n3915), .Q(n1265) );
  OAI2111 U5467 ( .A(n1266), .B(n3890), .C(n3864), .D(n3916), .Q(n3915) );
  AOI221 U5468 ( .A(n3866), .B(n3816), .C(n1323), .D(n3917), .Q(n3916) );
  XNR21 U5469 ( .A(n3968), .B(n3969), .Q(n3967) );
  INV3 U5470 ( .A(n3580), .Q(n1279) );
  INV3 U5471 ( .A(n3892), .Q(n1285) );
  INV3 U5472 ( .A(n4316), .Q(n1373) );
  INV3 U5473 ( .A(n3834), .Q(n1340) );
  AOI211 U5474 ( .A(n4265), .B(n3834), .C(n4086), .Q(n3453) );
  NOR21 U5475 ( .A(n3410), .B(n4069), .Q(n3859) );
  INV3 U5476 ( .A(n3862), .Q(n1238) );
  AOI221 U5477 ( .A(n1336), .B(n3861), .C(n1314), .D(n3664), .Q(n3860) );
  NAND22 U5478 ( .A(n4249), .B(n4250), .Q(n3862) );
  NAND22 U5479 ( .A(n4392), .B(n4393), .Q(n3814) );
  NAND22 U5480 ( .A(n4254), .B(n4255), .Q(n3861) );
  NAND22 U5481 ( .A(n3979), .B(n3980), .Q(n3612) );
  AOI221 U5482 ( .A(n1334), .B(n1254), .C(n1314), .D(n3837), .Q(n3980) );
  NAND22 U5483 ( .A(n4187), .B(n4188), .Q(n3982) );
  NAND22 U5484 ( .A(n4386), .B(n4387), .Q(n3575) );
  NAND22 U5485 ( .A(n4388), .B(n4389), .Q(n3815) );
  AOI221 U5486 ( .A(n6355), .B(n1456), .C(n1294), .D(n1453), .Q(n4388) );
  NAND22 U5487 ( .A(n4152), .B(n4153), .Q(n3396) );
  NAND22 U5488 ( .A(n4146), .B(n4147), .Q(n3800) );
  NAND22 U5489 ( .A(n4028), .B(n4029), .Q(n3931) );
  AOI221 U5490 ( .A(n1336), .B(n3395), .C(n1314), .D(n3800), .Q(n4029) );
  NAND22 U5491 ( .A(n4384), .B(n4385), .Q(n4065) );
  AOI221 U5492 ( .A(n1334), .B(n3814), .C(n1336), .D(n3921), .Q(n4384) );
  INV3 U5493 ( .A(n4006), .Q(n1353) );
  NAND22 U5494 ( .A(n3990), .B(n3991), .Q(n3705) );
  AOI221 U5495 ( .A(n1314), .B(n3861), .C(n1334), .D(n3664), .Q(n3991) );
  INV3 U5496 ( .A(n3766), .Q(n1348) );
  BUF2 U5497 ( .A(\execute/alu/sll_175/temp_int_SH[4] ), .Q(n6342) );
  AOI221 U5498 ( .A(n1314), .B(n1254), .C(n1336), .D(n3837), .Q(n3836) );
  AOI221 U5499 ( .A(n1336), .B(n3815), .C(n1314), .D(n3814), .Q(n3920) );
  NAND22 U5500 ( .A(n3941), .B(n3942), .Q(n3532) );
  NOR21 U5501 ( .A(n3919), .B(n3895), .Q(n4305) );
  INV3 U5502 ( .A(n3713), .Q(n1257) );
  INV3 U5503 ( .A(n6354), .Q(n6355) );
  INV3 U5504 ( .A(n3921), .Q(n1230) );
  NAND22 U5505 ( .A(n1174), .B(n6319), .Q(n6421) );
  NAND22 U5506 ( .A(n1163), .B(n6316), .Q(n6485) );
  NAND22 U5507 ( .A(n1174), .B(n6320), .Q(n6420) );
  NAND22 U5508 ( .A(n1163), .B(n6317), .Q(n6484) );
  NAND22 U5509 ( .A(n1174), .B(n6320), .Q(n1938) );
  NAND22 U5510 ( .A(n1163), .B(n6318), .Q(n2021) );
  NAND22 U5511 ( .A(n1173), .B(n6319), .Q(n6415) );
  NAND22 U5512 ( .A(n1172), .B(n6319), .Q(n6419) );
  NAND22 U5513 ( .A(n1166), .B(n6316), .Q(n6479) );
  NAND22 U5514 ( .A(n1165), .B(n6316), .Q(n6483) );
  NAND22 U5515 ( .A(n1173), .B(n6319), .Q(n6414) );
  NAND22 U5516 ( .A(n1172), .B(n6320), .Q(n6418) );
  NAND22 U5517 ( .A(n1166), .B(n6317), .Q(n6478) );
  NAND22 U5518 ( .A(n1165), .B(n6317), .Q(n6482) );
  NAND22 U5519 ( .A(n4086), .B(n1473), .Q(n3504) );
  NAND22 U5520 ( .A(n1173), .B(n6320), .Q(n1939) );
  NAND22 U5521 ( .A(n1172), .B(n6320), .Q(n1937) );
  NAND22 U5522 ( .A(n1166), .B(n6318), .Q(n2022) );
  NAND22 U5523 ( .A(n1165), .B(n6318), .Q(n2020) );
  INV3 U5524 ( .A(n6358), .Q(n1470) );
  NAND22 U5525 ( .A(n3606), .B(n3607), .Q(n3469) );
  INV3 U5526 ( .A(n3362), .Q(n1173) );
  INV3 U5527 ( .A(n2694), .Q(n1166) );
  NAND22 U5528 ( .A(n3703), .B(n3704), .Q(n3497) );
  NOR21 U5529 ( .A(n3362), .B(n6320), .Q(n6372) );
  INV3 U5530 ( .A(n3402), .Q(n6517) );
  BUF2 U5531 ( .A(n1943), .Q(n6407) );
  BUF2 U5532 ( .A(n1944), .Q(n6412) );
  BUF2 U5533 ( .A(n6404), .Q(n6406) );
  BUF2 U5534 ( .A(n6409), .Q(n6411) );
  BUF2 U5535 ( .A(n6404), .Q(n6405) );
  BUF2 U5536 ( .A(n6409), .Q(n6410) );
  BUF2 U5537 ( .A(n6468), .Q(n6470) );
  BUF2 U5538 ( .A(n6473), .Q(n6475) );
  BUF2 U5539 ( .A(n2026), .Q(n6471) );
  BUF2 U5540 ( .A(n2027), .Q(n6476) );
  BUF2 U5541 ( .A(n2026), .Q(n6472) );
  BUF2 U5542 ( .A(n2027), .Q(n6477) );
  BUF2 U5543 ( .A(n6468), .Q(n6469) );
  BUF2 U5544 ( .A(n6473), .Q(n6474) );
  BUF2 U5545 ( .A(n1943), .Q(n6408) );
  BUF2 U5546 ( .A(n1944), .Q(n6413) );
  INV3 U5547 ( .A(n6366), .Q(n6367) );
  INV3 U5548 ( .A(n6366), .Q(n6369) );
  INV3 U5549 ( .A(n6366), .Q(n6368) );
  INV3 U5550 ( .A(n6429), .Q(n6430) );
  INV3 U5551 ( .A(n6429), .Q(n6432) );
  INV3 U5552 ( .A(n6429), .Q(n6433) );
  INV3 U5553 ( .A(n6429), .Q(n6431) );
  INV3 U5554 ( .A(n6395), .Q(n6397) );
  INV3 U5555 ( .A(n6395), .Q(n6398) );
  INV3 U5556 ( .A(n6395), .Q(n6396) );
  INV3 U5557 ( .A(n6461), .Q(n6463) );
  INV3 U5558 ( .A(n6461), .Q(n6462) );
  INV3 U5559 ( .A(n6461), .Q(n6464) );
  INV3 U5560 ( .A(n3981), .Q(n1243) );
  BUF2 U5561 ( .A(n6384), .Q(n6387) );
  BUF2 U5562 ( .A(n6384), .Q(n6386) );
  BUF2 U5563 ( .A(n6447), .Q(n6449) );
  BUF2 U5564 ( .A(n6447), .Q(n6450) );
  INV3 U5565 ( .A(n6371), .Q(n6373) );
  NOR21 U5566 ( .A(n3362), .B(n6319), .Q(n6371) );
  NOR21 U5567 ( .A(n2694), .B(n6316), .Q(n2034) );
  INV3 U5568 ( .A(n6434), .Q(n6435) );
  NOR21 U5569 ( .A(n2694), .B(n6316), .Q(n6434) );
  INV3 U5570 ( .A(n6360), .Q(n6362) );
  INV3 U5571 ( .A(n6360), .Q(n6361) );
  INV3 U5572 ( .A(n6425), .Q(n6426) );
  INV3 U5573 ( .A(n6425), .Q(n6424) );
  INV3 U5574 ( .A(n6425), .Q(n6423) );
  INV3 U5575 ( .A(n6379), .Q(n6380) );
  INV3 U5576 ( .A(n6379), .Q(n6382) );
  INV3 U5577 ( .A(n6379), .Q(n6381) );
  INV3 U5578 ( .A(n6444), .Q(n6445) );
  INV3 U5579 ( .A(n6444), .Q(n6442) );
  INV3 U5580 ( .A(n6444), .Q(n6443) );
  INV3 U5581 ( .A(n4002), .Q(n1379) );
  BUF2 U5582 ( .A(n6385), .Q(n6389) );
  BUF2 U5583 ( .A(n6385), .Q(n6388) );
  BUF2 U5584 ( .A(n6448), .Q(n6452) );
  BUF2 U5585 ( .A(n2028), .Q(n6453) );
  BUF2 U5586 ( .A(n6448), .Q(n6451) );
  BUF2 U5587 ( .A(n1945), .Q(n6391) );
  BUF2 U5588 ( .A(n1945), .Q(n6390) );
  BUF2 U5589 ( .A(n2028), .Q(n6454) );
  NAND22 U5590 ( .A(n3739), .B(n3741), .Q(n3763) );
  INV3 U5591 ( .A(n6366), .Q(n6370) );
  INV3 U5592 ( .A(n3501), .Q(n1239) );
  INV3 U5593 ( .A(n6395), .Q(n6399) );
  INV3 U5594 ( .A(n6461), .Q(n6465) );
  INV3 U5595 ( .A(n6360), .Q(n6364) );
  INV3 U5596 ( .A(n6360), .Q(n6363) );
  INV3 U5597 ( .A(n6425), .Q(n6427) );
  INV3 U5598 ( .A(n6379), .Q(n6383) );
  INV3 U5599 ( .A(n6444), .Q(n6446) );
  INV3 U5600 ( .A(n4044), .Q(n1376) );
  INV3 U5601 ( .A(n3739), .Q(n1402) );
  INV3 U5602 ( .A(n6515), .Q(n6514) );
  INV3 U5603 ( .A(n3410), .Q(n1473) );
  INV3 U5604 ( .A(n3617), .Q(n1471) );
  BUF2 U5605 ( .A(n6726), .Q(n6722) );
  BUF2 U5606 ( .A(n6727), .Q(n6721) );
  BUF2 U5607 ( .A(n6727), .Q(n6720) );
  BUF2 U5608 ( .A(n6727), .Q(n6719) );
  BUF2 U5609 ( .A(n6727), .Q(n6718) );
  BUF2 U5610 ( .A(n6728), .Q(n6717) );
  BUF2 U5611 ( .A(n6728), .Q(n6716) );
  BUF2 U5612 ( .A(n6728), .Q(n6715) );
  BUF2 U5613 ( .A(n6728), .Q(n6714) );
  BUF2 U5614 ( .A(n6729), .Q(n6713) );
  BUF2 U5615 ( .A(n6729), .Q(n6712) );
  BUF2 U5616 ( .A(n6729), .Q(n6711) );
  BUF2 U5617 ( .A(n6729), .Q(n6710) );
  BUF2 U5618 ( .A(n6730), .Q(n6709) );
  BUF2 U5619 ( .A(n6730), .Q(n6708) );
  BUF2 U5620 ( .A(n6730), .Q(n6707) );
  BUF2 U5621 ( .A(n6730), .Q(n6706) );
  BUF2 U5622 ( .A(n6731), .Q(n6705) );
  BUF2 U5623 ( .A(n6731), .Q(n6704) );
  BUF2 U5624 ( .A(n6731), .Q(n6703) );
  BUF2 U5625 ( .A(n6731), .Q(n6702) );
  BUF2 U5626 ( .A(n6732), .Q(n6701) );
  BUF2 U5627 ( .A(n6732), .Q(n6700) );
  BUF2 U5628 ( .A(n6732), .Q(n6699) );
  BUF2 U5629 ( .A(n6732), .Q(n6698) );
  BUF2 U5630 ( .A(n6733), .Q(n6697) );
  BUF2 U5631 ( .A(n6733), .Q(n6696) );
  BUF2 U5632 ( .A(n6733), .Q(n6695) );
  BUF2 U5633 ( .A(n6733), .Q(n6694) );
  BUF2 U5634 ( .A(n6734), .Q(n6693) );
  BUF2 U5635 ( .A(n6734), .Q(n6692) );
  BUF2 U5636 ( .A(n6734), .Q(n6691) );
  BUF2 U5637 ( .A(n6734), .Q(n6690) );
  BUF2 U5638 ( .A(n6735), .Q(n6689) );
  BUF2 U5639 ( .A(n6735), .Q(n6688) );
  BUF2 U5640 ( .A(n6735), .Q(n6687) );
  BUF2 U5641 ( .A(n6735), .Q(n6686) );
  BUF2 U5642 ( .A(n6736), .Q(n6685) );
  BUF2 U5643 ( .A(n6736), .Q(n6684) );
  BUF2 U5644 ( .A(n6736), .Q(n6683) );
  BUF2 U5645 ( .A(n6736), .Q(n6682) );
  BUF2 U5646 ( .A(n6737), .Q(n6681) );
  BUF2 U5647 ( .A(n6737), .Q(n6680) );
  BUF2 U5648 ( .A(n6737), .Q(n6679) );
  BUF2 U5649 ( .A(n6737), .Q(n6678) );
  BUF2 U5650 ( .A(n6738), .Q(n6677) );
  BUF2 U5651 ( .A(n6738), .Q(n6676) );
  BUF2 U5652 ( .A(n6738), .Q(n6675) );
  BUF2 U5653 ( .A(n6738), .Q(n6674) );
  BUF2 U5654 ( .A(n6739), .Q(n6673) );
  BUF2 U5655 ( .A(n6739), .Q(n6672) );
  BUF2 U5656 ( .A(n6739), .Q(n6671) );
  BUF2 U5657 ( .A(n6739), .Q(n6670) );
  BUF2 U5658 ( .A(n6740), .Q(n6669) );
  BUF2 U5659 ( .A(n6740), .Q(n6668) );
  BUF2 U5660 ( .A(n6740), .Q(n6667) );
  BUF2 U5661 ( .A(n6740), .Q(n6666) );
  BUF2 U5662 ( .A(n6741), .Q(n6665) );
  BUF2 U5663 ( .A(n6741), .Q(n6664) );
  BUF2 U5664 ( .A(n6741), .Q(n6663) );
  BUF2 U5665 ( .A(n6741), .Q(n6662) );
  BUF2 U5666 ( .A(n6742), .Q(n6661) );
  BUF2 U5667 ( .A(n6742), .Q(n6660) );
  BUF2 U5668 ( .A(n6742), .Q(n6659) );
  BUF2 U5669 ( .A(n6742), .Q(n6658) );
  BUF2 U5670 ( .A(n6743), .Q(n6657) );
  BUF2 U5671 ( .A(n6743), .Q(n6656) );
  BUF2 U5672 ( .A(n6743), .Q(n6655) );
  BUF2 U5673 ( .A(n6743), .Q(n6654) );
  BUF2 U5674 ( .A(n6744), .Q(n6653) );
  BUF2 U5675 ( .A(n6744), .Q(n6652) );
  BUF2 U5676 ( .A(n6744), .Q(n6651) );
  BUF2 U5677 ( .A(n6744), .Q(n6650) );
  BUF2 U5678 ( .A(n6745), .Q(n6649) );
  BUF2 U5679 ( .A(n6745), .Q(n6648) );
  BUF2 U5680 ( .A(n6745), .Q(n6647) );
  BUF2 U5681 ( .A(n6745), .Q(n6646) );
  BUF2 U5682 ( .A(n6746), .Q(n6645) );
  BUF2 U5683 ( .A(n6746), .Q(n6644) );
  BUF2 U5684 ( .A(n6746), .Q(n6643) );
  BUF2 U5685 ( .A(n6746), .Q(n6642) );
  BUF2 U5686 ( .A(n6747), .Q(n6641) );
  BUF2 U5687 ( .A(n6747), .Q(n6640) );
  BUF2 U5688 ( .A(n6747), .Q(n6639) );
  BUF2 U5689 ( .A(n6747), .Q(n6638) );
  BUF2 U5690 ( .A(n6748), .Q(n6637) );
  BUF2 U5691 ( .A(n6748), .Q(n6636) );
  BUF2 U5692 ( .A(n6748), .Q(n6635) );
  BUF2 U5693 ( .A(n6748), .Q(n6634) );
  BUF2 U5694 ( .A(n6749), .Q(n6633) );
  BUF2 U5695 ( .A(n6749), .Q(n6632) );
  BUF2 U5696 ( .A(n6749), .Q(n6631) );
  BUF2 U5697 ( .A(n6749), .Q(n6630) );
  BUF2 U5698 ( .A(n6750), .Q(n6629) );
  BUF2 U5699 ( .A(n6750), .Q(n6628) );
  BUF2 U5700 ( .A(n6750), .Q(n6627) );
  BUF2 U5701 ( .A(n6750), .Q(n6626) );
  BUF2 U5702 ( .A(n6751), .Q(n6625) );
  BUF2 U5703 ( .A(n6751), .Q(n6624) );
  BUF2 U5704 ( .A(n6751), .Q(n6623) );
  BUF2 U5705 ( .A(n6751), .Q(n6622) );
  BUF2 U5706 ( .A(n6752), .Q(n6621) );
  BUF2 U5707 ( .A(n6752), .Q(n6620) );
  BUF2 U5708 ( .A(n6752), .Q(n6619) );
  BUF2 U5709 ( .A(n6752), .Q(n6618) );
  BUF2 U5710 ( .A(n6753), .Q(n6617) );
  BUF2 U5711 ( .A(n6753), .Q(n6616) );
  BUF2 U5712 ( .A(n6753), .Q(n6615) );
  BUF2 U5713 ( .A(n6753), .Q(n6614) );
  BUF2 U5714 ( .A(n6754), .Q(n6613) );
  BUF2 U5715 ( .A(n6754), .Q(n6612) );
  BUF2 U5716 ( .A(n6754), .Q(n6611) );
  BUF2 U5717 ( .A(n6754), .Q(n6610) );
  BUF2 U5718 ( .A(n6726), .Q(n6723) );
  BUF2 U5719 ( .A(n6726), .Q(n6724) );
  BUF2 U5720 ( .A(n6755), .Q(n6609) );
  BUF2 U5721 ( .A(n6755), .Q(n6608) );
  BUF2 U5722 ( .A(n6726), .Q(n6725) );
  INV3 U5723 ( .A(n3742), .Q(n1406) );
  NAND22 U5724 ( .A(n3827), .B(n1398), .Q(n3640) );
  XNR21 U5725 ( .A(n3911), .B(n6350), .Q(n3910) );
  NOR21 U5726 ( .A(n1447), .B(n1387), .Q(n4308) );
  INV3 U5727 ( .A(n4305), .Q(n1388) );
  NOR31 U5728 ( .A(n3846), .B(n1394), .C(n1390), .Q(n3805) );
  NAND31 U5729 ( .A(n1385), .B(n1383), .C(n1381), .Q(n4475) );
  NAND31 U5730 ( .A(n1408), .B(n1404), .C(n1405), .Q(n4474) );
  NAND22 U5731 ( .A(n4240), .B(n1351), .Q(n4055) );
  INV3 U5732 ( .A(n6331), .Q(n6333) );
  INV3 U5733 ( .A(n6328), .Q(n6330) );
  NAND22 U5734 ( .A(n3668), .B(n3669), .Q(n3643) );
  XOR21 U5735 ( .A(n6321), .B(n1439), .Q(n6261) );
  BUF2 U5736 ( .A(\instruction_decode/reg_MAPP/n1245 ), .Q(n6763) );
  BUF2 U5737 ( .A(\instruction_decode/reg_MAPP/n1245 ), .Q(n6764) );
  BUF2 U5738 ( .A(\instruction_decode/reg_MAPP/n1245 ), .Q(n6765) );
  BUF2 U5739 ( .A(\instruction_decode/reg_MAPP/n1245 ), .Q(n6766) );
  BUF2 U5740 ( .A(\instruction_decode/reg_MAPP/n1272 ), .Q(n6899) );
  BUF2 U5741 ( .A(\instruction_decode/reg_MAPP/n1272 ), .Q(n6900) );
  BUF2 U5742 ( .A(\instruction_decode/reg_MAPP/n1272 ), .Q(n6901) );
  BUF2 U5743 ( .A(\instruction_decode/reg_MAPP/n1261 ), .Q(n6843) );
  BUF2 U5744 ( .A(\instruction_decode/reg_MAPP/n1261 ), .Q(n6844) );
  BUF2 U5745 ( .A(\instruction_decode/reg_MAPP/n1261 ), .Q(n6845) );
  BUF2 U5746 ( .A(\instruction_decode/reg_MAPP/n1261 ), .Q(n6846) );
  BUF2 U5747 ( .A(\instruction_decode/reg_MAPP/n1253 ), .Q(n6803) );
  BUF2 U5748 ( .A(\instruction_decode/reg_MAPP/n1253 ), .Q(n6804) );
  BUF2 U5749 ( .A(\instruction_decode/reg_MAPP/n1253 ), .Q(n6805) );
  BUF2 U5750 ( .A(\instruction_decode/reg_MAPP/n1253 ), .Q(n6806) );
  BUF2 U5751 ( .A(\instruction_decode/reg_MAPP/n1272 ), .Q(n6898) );
  BUF2 U5752 ( .A(\instruction_decode/reg_MAPP/n1245 ), .Q(n6767) );
  BUF2 U5753 ( .A(\instruction_decode/reg_MAPP/n1261 ), .Q(n6847) );
  BUF2 U5754 ( .A(\instruction_decode/reg_MAPP/n1253 ), .Q(n6807) );
  BUF2 U5755 ( .A(\instruction_decode/reg_MAPP/n1272 ), .Q(n6902) );
  AOI211 U5756 ( .A(n3644), .B(n1353), .C(n3645), .Q(n3618) );
  XNR21 U5757 ( .A(n3755), .B(n3627), .Q(n3737) );
  XNR21 U5758 ( .A(n3716), .B(n6350), .Q(n3670) );
  NAND22 U5759 ( .A(n1413), .B(n1356), .Q(n4350) );
  XNR21 U5760 ( .A(n3793), .B(n3627), .Q(n3806) );
  NAND22 U5761 ( .A(n1413), .B(n4394), .Q(n4401) );
  NAND22 U5762 ( .A(n3825), .B(n1401), .Q(n3641) );
  OAI2111 U5763 ( .A(n3778), .B(n3779), .C(n6352), .D(n3780), .Q(n3776) );
  NAND22 U5764 ( .A(n6513), .B(n1455), .Q(n3779) );
  XNR21 U5765 ( .A(n4077), .B(n4078), .Q(n4076) );
  NOR40 U5766 ( .A(n3853), .B(n3854), .C(n3855), .D(n3856), .Q(n3852) );
  NAND22 U5767 ( .A(n3970), .B(n1387), .Q(n3912) );
  NAND22 U5768 ( .A(n1259), .B(n1310), .Q(n4256) );
  NAND41 U5769 ( .A(n4030), .B(n4031), .C(n4032), .D(n4033), .Q(
        \execute/old_res [16]) );
  NAND22 U5770 ( .A(n6236), .B(n4065), .Q(n4031) );
  NAND41 U5771 ( .A(n3520), .B(n3521), .C(n3522), .D(n3523), .Q(
        \execute/old_res [5]) );
  NOR40 U5772 ( .A(n4158), .B(n4159), .C(n4160), .D(n4161), .Q(n4157) );
  NOR40 U5773 ( .A(n3524), .B(n1249), .C(n1221), .D(n3525), .Q(n3523) );
  INV3 U5774 ( .A(n3531), .Q(n1249) );
  NOR40 U5775 ( .A(n4117), .B(n4118), .C(n4119), .D(n4120), .Q(n4116) );
  AOI2111 U5776 ( .A(n1316), .B(n3664), .C(n4103), .D(n4104), .Q(n4095) );
  INV3 U5777 ( .A(n4082), .Q(n1316) );
  NAND22 U5778 ( .A(n3726), .B(n1409), .Q(n3672) );
  AOI221 U5779 ( .A(\execute/alu/sll_175/ML_int[5][23] ), .B(n1353), .C(n6236), 
        .D(n3486), .Q(n3835) );
  INV3 U5780 ( .A(n4102), .Q(n1324) );
  AOI221 U5781 ( .A(\execute/alu/sll_175/ML_int[4][14] ), .B(n1341), .C(n4101), 
        .D(n6515), .Q(n4100) );
  NAND22 U5782 ( .A(n3670), .B(n1410), .Q(n3668) );
  NAND31 U5783 ( .A(n4010), .B(n4011), .C(n4012), .Q(\execute/old_res [17]) );
  AOI2111 U5784 ( .A(n1443), .B(n4013), .C(n4014), .D(n4015), .Q(n4012) );
  AOI221 U5785 ( .A(n3859), .B(n3954), .C(\execute/alu/sll_175/ML_int[5][17] ), 
        .D(n1353), .Q(n4011) );
  AOI221 U5786 ( .A(n1218), .B(n3507), .C(n3687), .D(n6513), .Q(n3686) );
  XNR21 U5787 ( .A(n3590), .B(n3688), .Q(n3687) );
  NOR21 U5788 ( .A(n3825), .B(n1401), .Q(n3642) );
  XNR21 U5789 ( .A(n4109), .B(n4080), .Q(n4108) );
  NAND22 U5790 ( .A(n1375), .B(n4057), .Q(n4109) );
  INV3 U5791 ( .A(n3631), .Q(n1412) );
  INV3 U5792 ( .A(n3971), .Q(n1386) );
  NAND22 U5793 ( .A(n4070), .B(n4071), .Q(\execute/old_res [15]) );
  NOR40 U5794 ( .A(n1241), .B(n4088), .C(n4089), .D(n4090), .Q(n4070) );
  NOR40 U5795 ( .A(n4072), .B(n4073), .C(n4074), .D(n4075), .Q(n4071) );
  BUF2 U5796 ( .A(\instruction_decode/reg_MAPP/n1275 ), .Q(n6913) );
  BUF2 U5797 ( .A(\instruction_decode/reg_MAPP/n1275 ), .Q(n6914) );
  BUF2 U5798 ( .A(\instruction_decode/reg_MAPP/n1275 ), .Q(n6915) );
  BUF2 U5799 ( .A(\instruction_decode/reg_MAPP/n1275 ), .Q(n6916) );
  BUF2 U5800 ( .A(\instruction_decode/reg_MAPP/n1269 ), .Q(n6883) );
  BUF2 U5801 ( .A(\instruction_decode/reg_MAPP/n1269 ), .Q(n6884) );
  BUF2 U5802 ( .A(\instruction_decode/reg_MAPP/n1269 ), .Q(n6885) );
  BUF2 U5803 ( .A(\instruction_decode/reg_MAPP/n1269 ), .Q(n6886) );
  BUF2 U5804 ( .A(\instruction_decode/reg_MAPP/n1273 ), .Q(n6903) );
  BUF2 U5805 ( .A(\instruction_decode/reg_MAPP/n1273 ), .Q(n6904) );
  BUF2 U5806 ( .A(\instruction_decode/reg_MAPP/n1273 ), .Q(n6905) );
  BUF2 U5807 ( .A(\instruction_decode/reg_MAPP/n1273 ), .Q(n6906) );
  BUF2 U5808 ( .A(\instruction_decode/reg_MAPP/n1248 ), .Q(n6778) );
  BUF2 U5809 ( .A(\instruction_decode/reg_MAPP/n1248 ), .Q(n6779) );
  BUF2 U5810 ( .A(\instruction_decode/reg_MAPP/n1248 ), .Q(n6780) );
  BUF2 U5811 ( .A(\instruction_decode/reg_MAPP/n1248 ), .Q(n6781) );
  BUF2 U5812 ( .A(\instruction_decode/reg_MAPP/n1264 ), .Q(n6858) );
  BUF2 U5813 ( .A(\instruction_decode/reg_MAPP/n1264 ), .Q(n6859) );
  BUF2 U5814 ( .A(\instruction_decode/reg_MAPP/n1264 ), .Q(n6860) );
  BUF2 U5815 ( .A(\instruction_decode/reg_MAPP/n1264 ), .Q(n6861) );
  BUF2 U5816 ( .A(\instruction_decode/reg_MAPP/n1256 ), .Q(n6818) );
  BUF2 U5817 ( .A(\instruction_decode/reg_MAPP/n1256 ), .Q(n6819) );
  BUF2 U5818 ( .A(\instruction_decode/reg_MAPP/n1256 ), .Q(n6820) );
  BUF2 U5819 ( .A(\instruction_decode/reg_MAPP/n1256 ), .Q(n6821) );
  BUF2 U5820 ( .A(\instruction_decode/reg_MAPP/n1250 ), .Q(n6788) );
  BUF2 U5821 ( .A(\instruction_decode/reg_MAPP/n1250 ), .Q(n6789) );
  BUF2 U5822 ( .A(\instruction_decode/reg_MAPP/n1250 ), .Q(n6790) );
  BUF2 U5823 ( .A(\instruction_decode/reg_MAPP/n1250 ), .Q(n6791) );
  BUF2 U5824 ( .A(\instruction_decode/reg_MAPP/n1266 ), .Q(n6868) );
  BUF2 U5825 ( .A(\instruction_decode/reg_MAPP/n1266 ), .Q(n6869) );
  BUF2 U5826 ( .A(\instruction_decode/reg_MAPP/n1266 ), .Q(n6870) );
  BUF2 U5827 ( .A(\instruction_decode/reg_MAPP/n1266 ), .Q(n6871) );
  BUF2 U5828 ( .A(\instruction_decode/reg_MAPP/n1258 ), .Q(n6828) );
  BUF2 U5829 ( .A(\instruction_decode/reg_MAPP/n1258 ), .Q(n6829) );
  BUF2 U5830 ( .A(\instruction_decode/reg_MAPP/n1258 ), .Q(n6830) );
  BUF2 U5831 ( .A(\instruction_decode/reg_MAPP/n1258 ), .Q(n6831) );
  BUF2 U5832 ( .A(\instruction_decode/reg_MAPP/n1246 ), .Q(n6768) );
  BUF2 U5833 ( .A(\instruction_decode/reg_MAPP/n1246 ), .Q(n6769) );
  BUF2 U5834 ( .A(\instruction_decode/reg_MAPP/n1246 ), .Q(n6770) );
  BUF2 U5835 ( .A(\instruction_decode/reg_MAPP/n1246 ), .Q(n6771) );
  BUF2 U5836 ( .A(\instruction_decode/reg_MAPP/n1262 ), .Q(n6848) );
  BUF2 U5837 ( .A(\instruction_decode/reg_MAPP/n1262 ), .Q(n6849) );
  BUF2 U5838 ( .A(\instruction_decode/reg_MAPP/n1262 ), .Q(n6850) );
  BUF2 U5839 ( .A(\instruction_decode/reg_MAPP/n1262 ), .Q(n6851) );
  BUF2 U5840 ( .A(\instruction_decode/reg_MAPP/n1254 ), .Q(n6808) );
  BUF2 U5841 ( .A(\instruction_decode/reg_MAPP/n1254 ), .Q(n6809) );
  BUF2 U5842 ( .A(\instruction_decode/reg_MAPP/n1254 ), .Q(n6810) );
  BUF2 U5843 ( .A(\instruction_decode/reg_MAPP/n1254 ), .Q(n6811) );
  BUF2 U5844 ( .A(\instruction_decode/reg_MAPP/n1275 ), .Q(n6917) );
  BUF2 U5845 ( .A(\instruction_decode/reg_MAPP/n1269 ), .Q(n6887) );
  BUF2 U5846 ( .A(\instruction_decode/reg_MAPP/n1273 ), .Q(n6907) );
  BUF2 U5847 ( .A(\instruction_decode/reg_MAPP/n1248 ), .Q(n6782) );
  BUF2 U5848 ( .A(\instruction_decode/reg_MAPP/n1264 ), .Q(n6862) );
  BUF2 U5849 ( .A(\instruction_decode/reg_MAPP/n1256 ), .Q(n6822) );
  BUF2 U5850 ( .A(\instruction_decode/reg_MAPP/n1250 ), .Q(n6792) );
  BUF2 U5851 ( .A(\instruction_decode/reg_MAPP/n1266 ), .Q(n6872) );
  BUF2 U5852 ( .A(\instruction_decode/reg_MAPP/n1258 ), .Q(n6832) );
  BUF2 U5853 ( .A(\instruction_decode/reg_MAPP/n1246 ), .Q(n6772) );
  BUF2 U5854 ( .A(\instruction_decode/reg_MAPP/n1262 ), .Q(n6852) );
  BUF2 U5855 ( .A(\instruction_decode/reg_MAPP/n1254 ), .Q(n6812) );
  AOI221 U5856 ( .A(\execute/alu/sll_175/ML_int[5][24] ), .B(n1353), .C(n6236), 
        .D(n1229), .Q(n3813) );
  INV3 U5857 ( .A(n3446), .Q(n1229) );
  NAND31 U5858 ( .A(n4068), .B(n1342), .C(n4067), .Q(n3569) );
  AOI211 U5859 ( .A(n6515), .B(n1310), .C(n3952), .Q(n3951) );
  NOR21 U5860 ( .A(n1330), .B(n4270), .Q(n3866) );
  NAND22 U5861 ( .A(n5821), .B(n4400), .Q(n3611) );
  NAND22 U5862 ( .A(n4087), .B(n6234), .Q(n4069) );
  NAND22 U5863 ( .A(n4355), .B(n4270), .Q(n3863) );
  OAI2111 U5864 ( .A(n4021), .B(n3407), .C(n4022), .D(n3766), .Q(n4014) );
  NAND22 U5865 ( .A(n5821), .B(n1290), .Q(n3610) );
  AOI221 U5866 ( .A(n1325), .B(n3571), .C(n1349), .D(n4065), .Q(n4383) );
  NOR21 U5867 ( .A(n4350), .B(n4087), .Q(n4265) );
  NAND41 U5868 ( .A(n3492), .B(n3493), .C(n3494), .D(n3495), .Q(n3491) );
  NOR21 U5869 ( .A(n4400), .B(n5821), .Q(n3615) );
  NOR40 U5870 ( .A(n3984), .B(n3985), .C(n3986), .D(n3987), .Q(n3983) );
  NOR21 U5871 ( .A(n1413), .B(n1357), .Q(n4458) );
  INV3 U5872 ( .A(n4480), .Q(n1357) );
  NAND41 U5873 ( .A(n4481), .B(n4482), .C(n4483), .D(n4484), .Q(n4480) );
  NOR40 U5874 ( .A(n4500), .B(n1381), .C(n1395), .D(n1387), .Q(n4483) );
  INV3 U5875 ( .A(n3571), .Q(n1261) );
  NAND22 U5876 ( .A(n4271), .B(n4272), .Q(n3513) );
  INV3 U5877 ( .A(n3481), .Q(n1275) );
  INV3 U5878 ( .A(n3394), .Q(n1250) );
  NAND41 U5879 ( .A(n3576), .B(n3577), .C(n3578), .D(n3579), .Q(
        \execute/old_res [3]) );
  NAND41 U5880 ( .A(n4218), .B(n4219), .C(n4220), .D(n4221), .Q(
        \execute/old_res [10]) );
  NAND22 U5881 ( .A(n6512), .B(n1428), .Q(n4219) );
  NAND22 U5882 ( .A(n4000), .B(n1379), .Q(n4019) );
  NAND41 U5883 ( .A(n4260), .B(n3453), .C(n4261), .D(n1273), .Q(n4259) );
  NOR21 U5884 ( .A(n4270), .B(n4355), .Q(n3994) );
  NAND22 U5885 ( .A(n4358), .B(n4359), .Q(n3917) );
  AOI221 U5886 ( .A(n6516), .B(n1443), .C(n6515), .D(n4018), .Q(n4017) );
  NAND31 U5887 ( .A(n1444), .B(n4019), .C(n6513), .Q(n4016) );
  INV3 U5888 ( .A(n3511), .Q(n1300) );
  INV3 U5889 ( .A(n3505), .Q(n1219) );
  INV3 U5890 ( .A(n3931), .Q(n1246) );
  AOI221 U5891 ( .A(n1331), .B(n4178), .C(n1328), .D(n3574), .Q(n4345) );
  INV3 U5892 ( .A(n4066), .Q(n1262) );
  NOR40 U5893 ( .A(n3450), .B(n3451), .C(n1339), .D(n3452), .Q(n3448) );
  NAND22 U5894 ( .A(n4192), .B(n4193), .Q(n3485) );
  NAND22 U5895 ( .A(n4123), .B(n4124), .Q(n3892) );
  INV3 U5896 ( .A(n3480), .Q(n1276) );
  INV3 U5897 ( .A(n3953), .Q(n1282) );
  INV3 U5898 ( .A(n3509), .Q(n1301) );
  AOI2111 U5899 ( .A(n1336), .B(n3497), .C(n3699), .D(n3700), .Q(n3695) );
  INV3 U5900 ( .A(n3563), .Q(n1352) );
  XNR21 U5901 ( .A(n3622), .B(n1413), .Q(n3625) );
  NAND22 U5902 ( .A(n3483), .B(n3453), .Q(n3478) );
  AOI211 U5903 ( .A(n1302), .B(n1423), .C(n1356), .Q(n3517) );
  NAND31 U5904 ( .A(n3922), .B(n3923), .C(n3924), .Q(\execute/old_res [1]) );
  AOI211 U5905 ( .A(n1325), .B(n3530), .C(n1282), .Q(n3922) );
  INV3 U5906 ( .A(n4355), .Q(n1330) );
  NAND22 U5907 ( .A(n3449), .B(n3421), .Q(n4325) );
  NOR21 U5908 ( .A(n4101), .B(n1378), .Q(n4316) );
  INV3 U5909 ( .A(n4400), .Q(n1290) );
  INV3 U5910 ( .A(n4237), .Q(n1297) );
  INV3 U5911 ( .A(n3484), .Q(n1277) );
  INV3 U5912 ( .A(n4178), .Q(n1268) );
  INV3 U5913 ( .A(n3545), .Q(n1284) );
  INV3 U5914 ( .A(n3574), .Q(n1269) );
  INV3 U5915 ( .A(n3536), .Q(n1287) );
  BUF2 U5916 ( .A(\instruction_decode/reg_MAPP/n1271 ), .Q(n6893) );
  BUF2 U5917 ( .A(\instruction_decode/reg_MAPP/n1271 ), .Q(n6894) );
  BUF2 U5918 ( .A(\instruction_decode/reg_MAPP/n1271 ), .Q(n6895) );
  BUF2 U5919 ( .A(\instruction_decode/reg_MAPP/n1271 ), .Q(n6896) );
  BUF2 U5920 ( .A(\instruction_decode/reg_MAPP/n1252 ), .Q(n6798) );
  BUF2 U5921 ( .A(\instruction_decode/reg_MAPP/n1252 ), .Q(n6799) );
  BUF2 U5922 ( .A(\instruction_decode/reg_MAPP/n1252 ), .Q(n6800) );
  BUF2 U5923 ( .A(\instruction_decode/reg_MAPP/n1252 ), .Q(n6801) );
  BUF2 U5924 ( .A(\instruction_decode/reg_MAPP/n1268 ), .Q(n6878) );
  BUF2 U5925 ( .A(\instruction_decode/reg_MAPP/n1268 ), .Q(n6879) );
  BUF2 U5926 ( .A(\instruction_decode/reg_MAPP/n1268 ), .Q(n6880) );
  BUF2 U5927 ( .A(\instruction_decode/reg_MAPP/n1268 ), .Q(n6881) );
  BUF2 U5928 ( .A(\instruction_decode/reg_MAPP/n1260 ), .Q(n6839) );
  BUF2 U5929 ( .A(\instruction_decode/reg_MAPP/n1260 ), .Q(n6840) );
  BUF2 U5930 ( .A(\instruction_decode/reg_MAPP/n1260 ), .Q(n6841) );
  BUF2 U5931 ( .A(\instruction_decode/reg_MAPP/n1260 ), .Q(n6838) );
  BUF2 U5932 ( .A(\instruction_decode/reg_MAPP/n1255 ), .Q(n6813) );
  BUF2 U5933 ( .A(\instruction_decode/reg_MAPP/n1255 ), .Q(n6814) );
  BUF2 U5934 ( .A(\instruction_decode/reg_MAPP/n1255 ), .Q(n6815) );
  BUF2 U5935 ( .A(\instruction_decode/reg_MAPP/n1255 ), .Q(n6816) );
  BUF2 U5936 ( .A(\instruction_decode/reg_MAPP/n1259 ), .Q(n6835) );
  BUF2 U5937 ( .A(\instruction_decode/reg_MAPP/n1259 ), .Q(n6836) );
  BUF2 U5938 ( .A(\instruction_decode/reg_MAPP/n1257 ), .Q(n6824) );
  BUF2 U5939 ( .A(\instruction_decode/reg_MAPP/n1257 ), .Q(n6825) );
  BUF2 U5940 ( .A(\instruction_decode/reg_MAPP/n1257 ), .Q(n6826) );
  BUF2 U5941 ( .A(\instruction_decode/reg_MAPP/n1259 ), .Q(n6834) );
  BUF2 U5942 ( .A(\instruction_decode/reg_MAPP/n1259 ), .Q(n6833) );
  BUF2 U5943 ( .A(\instruction_decode/reg_MAPP/n1257 ), .Q(n6823) );
  BUF2 U5944 ( .A(\instruction_decode/reg_MAPP/n1267 ), .Q(n6873) );
  BUF2 U5945 ( .A(\instruction_decode/reg_MAPP/n1267 ), .Q(n6874) );
  BUF2 U5946 ( .A(\instruction_decode/reg_MAPP/n1267 ), .Q(n6875) );
  BUF2 U5947 ( .A(\instruction_decode/reg_MAPP/n1267 ), .Q(n6876) );
  BUF2 U5948 ( .A(\instruction_decode/reg_MAPP/n1265 ), .Q(n6863) );
  BUF2 U5949 ( .A(\instruction_decode/reg_MAPP/n1265 ), .Q(n6864) );
  BUF2 U5950 ( .A(\instruction_decode/reg_MAPP/n1265 ), .Q(n6865) );
  BUF2 U5951 ( .A(\instruction_decode/reg_MAPP/n1265 ), .Q(n6866) );
  BUF2 U5952 ( .A(\instruction_decode/reg_MAPP/n1263 ), .Q(n6853) );
  BUF2 U5953 ( .A(\instruction_decode/reg_MAPP/n1263 ), .Q(n6854) );
  BUF2 U5954 ( .A(\instruction_decode/reg_MAPP/n1263 ), .Q(n6855) );
  BUF2 U5955 ( .A(\instruction_decode/reg_MAPP/n1263 ), .Q(n6856) );
  BUF2 U5956 ( .A(\instruction_decode/reg_MAPP/n1251 ), .Q(n6793) );
  BUF2 U5957 ( .A(\instruction_decode/reg_MAPP/n1251 ), .Q(n6794) );
  BUF2 U5958 ( .A(\instruction_decode/reg_MAPP/n1251 ), .Q(n6795) );
  BUF2 U5959 ( .A(\instruction_decode/reg_MAPP/n1251 ), .Q(n6796) );
  BUF2 U5960 ( .A(\instruction_decode/reg_MAPP/n1249 ), .Q(n6783) );
  BUF2 U5961 ( .A(\instruction_decode/reg_MAPP/n1249 ), .Q(n6784) );
  BUF2 U5962 ( .A(\instruction_decode/reg_MAPP/n1249 ), .Q(n6785) );
  BUF2 U5963 ( .A(\instruction_decode/reg_MAPP/n1249 ), .Q(n6786) );
  BUF2 U5964 ( .A(\instruction_decode/reg_MAPP/n1247 ), .Q(n6773) );
  BUF2 U5965 ( .A(\instruction_decode/reg_MAPP/n1247 ), .Q(n6774) );
  BUF2 U5966 ( .A(\instruction_decode/reg_MAPP/n1247 ), .Q(n6775) );
  BUF2 U5967 ( .A(\instruction_decode/reg_MAPP/n1247 ), .Q(n6776) );
  BUF2 U5968 ( .A(\instruction_decode/reg_MAPP/n1274 ), .Q(n6908) );
  BUF2 U5969 ( .A(\instruction_decode/reg_MAPP/n1274 ), .Q(n6909) );
  BUF2 U5970 ( .A(\instruction_decode/reg_MAPP/n1274 ), .Q(n6910) );
  BUF2 U5971 ( .A(\instruction_decode/reg_MAPP/n1274 ), .Q(n6911) );
  BUF2 U5972 ( .A(\instruction_decode/reg_MAPP/n1270 ), .Q(n6889) );
  BUF2 U5973 ( .A(\instruction_decode/reg_MAPP/n1270 ), .Q(n6890) );
  BUF2 U5974 ( .A(\instruction_decode/reg_MAPP/n1270 ), .Q(n6891) );
  BUF2 U5975 ( .A(\instruction_decode/reg_MAPP/n1276 ), .Q(n6918) );
  BUF2 U5976 ( .A(\instruction_decode/reg_MAPP/n1276 ), .Q(n6919) );
  BUF2 U5977 ( .A(\instruction_decode/reg_MAPP/n1276 ), .Q(n6920) );
  BUF2 U5978 ( .A(\instruction_decode/reg_MAPP/n1276 ), .Q(n6921) );
  BUF2 U5979 ( .A(\instruction_decode/reg_MAPP/n1270 ), .Q(n6888) );
  INV3 U5980 ( .A(n3518), .Q(n1272) );
  INV3 U5981 ( .A(n4216), .Q(n1296) );
  BUF2 U5982 ( .A(\instruction_decode/reg_MAPP/n1271 ), .Q(n6897) );
  BUF2 U5983 ( .A(\instruction_decode/reg_MAPP/n1252 ), .Q(n6802) );
  BUF2 U5984 ( .A(\instruction_decode/reg_MAPP/n1268 ), .Q(n6882) );
  BUF2 U5985 ( .A(\instruction_decode/reg_MAPP/n1260 ), .Q(n6842) );
  BUF2 U5986 ( .A(\instruction_decode/reg_MAPP/n1255 ), .Q(n6817) );
  BUF2 U5987 ( .A(\instruction_decode/reg_MAPP/n1259 ), .Q(n6837) );
  BUF2 U5988 ( .A(\instruction_decode/reg_MAPP/n1257 ), .Q(n6827) );
  BUF2 U5989 ( .A(\instruction_decode/reg_MAPP/n1267 ), .Q(n6877) );
  BUF2 U5990 ( .A(\instruction_decode/reg_MAPP/n1265 ), .Q(n6867) );
  BUF2 U5991 ( .A(\instruction_decode/reg_MAPP/n1263 ), .Q(n6857) );
  BUF2 U5992 ( .A(\instruction_decode/reg_MAPP/n1251 ), .Q(n6797) );
  BUF2 U5993 ( .A(\instruction_decode/reg_MAPP/n1249 ), .Q(n6787) );
  BUF2 U5994 ( .A(\instruction_decode/reg_MAPP/n1247 ), .Q(n6777) );
  BUF2 U5995 ( .A(\instruction_decode/reg_MAPP/n1274 ), .Q(n6912) );
  BUF2 U5996 ( .A(\instruction_decode/reg_MAPP/n1270 ), .Q(n6892) );
  BUF2 U5997 ( .A(\instruction_decode/reg_MAPP/n1276 ), .Q(n6922) );
  INV3 U5998 ( .A(n4131), .Q(n1294) );
  OAI2111 U5999 ( .A(n3407), .B(n3432), .C(n3433), .D(n3434), .Q(n3428) );
  INV3 U6000 ( .A(n3572), .Q(n1228) );
  NAND31 U6001 ( .A(n6513), .B(n6250), .C(n3474), .Q(n3511) );
  NAND22 U6002 ( .A(n4067), .B(n4068), .Q(n4006) );
  INV3 U6003 ( .A(inst_out[20]), .Q(n6317) );
  INV3 U6004 ( .A(n3390), .Q(n1349) );
  INV3 U6005 ( .A(n3500), .Q(n1235) );
  NAND22 U6006 ( .A(n4390), .B(n4391), .Q(n3921) );
  NAND22 U6007 ( .A(n4148), .B(n4149), .Q(n3395) );
  AOI221 U6008 ( .A(n6516), .B(n6222), .C(n6515), .D(n4039), .Q(n4038) );
  NOR21 U6009 ( .A(n6222), .B(n6357), .Q(n4043) );
  INV3 U6010 ( .A(n3999), .Q(n1445) );
  AOI221 U6011 ( .A(n6236), .B(n3933), .C(n3934), .D(n6513), .Q(n3932) );
  XNR21 U6012 ( .A(n3693), .B(n3935), .Q(n3934) );
  OAI2111 U6013 ( .A(n1251), .B(n3605), .C(n1252), .D(n3940), .Q(n3933) );
  NAND22 U6014 ( .A(n4228), .B(n4229), .Q(n3501) );
  NAND22 U6015 ( .A(n3602), .B(n1458), .Q(n4209) );
  INV3 U6016 ( .A(n3972), .Q(n1447) );
  AOI221 U6017 ( .A(n1336), .B(n3532), .C(n1334), .D(n3394), .Q(n3940) );
  INV3 U6018 ( .A(n3911), .Q(n1448) );
  NAND31 U6019 ( .A(n6352), .B(n3511), .C(n3514), .Q(n3512) );
  AOI221 U6020 ( .A(n6516), .B(n6193), .C(n6515), .D(n6348), .Q(n3514) );
  BUF2 U6021 ( .A(n3602), .Q(n6356) );
  NOR21 U6022 ( .A(n1449), .B(n1395), .Q(n3895) );
  NOR21 U6023 ( .A(n1448), .B(n1393), .Q(n3919) );
  INV3 U6024 ( .A(n3407), .Q(n6513) );
  NOR21 U6025 ( .A(n1259), .B(n1310), .Q(n6353) );
  INV3 U6026 ( .A(n3603), .Q(n6354) );
  NOR21 U6027 ( .A(n1259), .B(n1310), .Q(n3603) );
  INV3 U6028 ( .A(n3427), .Q(n1234) );
  INV3 U6029 ( .A(n3502), .Q(n1237) );
  INV3 U6030 ( .A(n3460), .Q(n1242) );
  INV3 U6031 ( .A(n3423), .Q(n1251) );
  INV3 U6032 ( .A(n3369), .Q(n1170) );
  NOR21 U6033 ( .A(n3365), .B(n6320), .Q(n3369) );
  INV3 U6034 ( .A(n2701), .Q(n1162) );
  NOR21 U6035 ( .A(n2697), .B(n6318), .Q(n2701) );
  NAND22 U6036 ( .A(n3359), .B(n3372), .Q(n3362) );
  NAND22 U6037 ( .A(n2691), .B(n2704), .Q(n2694) );
  NAND22 U6038 ( .A(n1161), .B(n6492), .Q(n6458) );
  NAND22 U6039 ( .A(n1161), .B(n6492), .Q(n6457) );
  NAND22 U6040 ( .A(n1171), .B(n6498), .Q(n6401) );
  NAND22 U6041 ( .A(n1171), .B(n6498), .Q(n6400) );
  NAND22 U6042 ( .A(n1175), .B(n6319), .Q(n6417) );
  NAND22 U6043 ( .A(n1164), .B(n6316), .Q(n6481) );
  NAND22 U6044 ( .A(n1161), .B(n6316), .Q(n6467) );
  NAND22 U6045 ( .A(n1169), .B(n6320), .Q(n1941) );
  NAND22 U6046 ( .A(n1175), .B(n6320), .Q(n6416) );
  NAND22 U6047 ( .A(n1169), .B(n6320), .Q(n6402) );
  NAND22 U6048 ( .A(n1164), .B(n6317), .Q(n6480) );
  NAND22 U6049 ( .A(n1161), .B(n6317), .Q(n6466) );
  NAND22 U6050 ( .A(n1171), .B(n6498), .Q(n1948) );
  NAND22 U6051 ( .A(n1161), .B(n6492), .Q(n2033) );
  NOR21 U6052 ( .A(n4395), .B(n1478), .Q(n3402) );
  NAND22 U6053 ( .A(n1169), .B(n6319), .Q(n6403) );
  NAND22 U6054 ( .A(n1175), .B(n6320), .Q(n1940) );
  NAND22 U6055 ( .A(n1164), .B(n6318), .Q(n2023) );
  NAND22 U6056 ( .A(n1161), .B(n6318), .Q(n2024) );
  NAND22 U6057 ( .A(n1175), .B(n6498), .Q(n6393) );
  NAND22 U6058 ( .A(n1175), .B(n6498), .Q(n6392) );
  NAND22 U6059 ( .A(n1164), .B(n6492), .Q(n6456) );
  NAND22 U6060 ( .A(n1164), .B(n6492), .Q(n6455) );
  INV3 U6061 ( .A(n6496), .Q(n6316) );
  INV3 U6062 ( .A(n6497), .Q(n6319) );
  AOI211 U6063 ( .A(n6515), .B(n1344), .C(n6512), .Q(n3559) );
  NAND22 U6064 ( .A(n1175), .B(n6498), .Q(n1949) );
  NAND22 U6065 ( .A(n1164), .B(n6492), .Q(n2032) );
  INV3 U6066 ( .A(n6497), .Q(n6320) );
  INV3 U6067 ( .A(n6496), .Q(n6318) );
  INV3 U6068 ( .A(n4372), .Q(n1336) );
  OAI2111 U6069 ( .A(n3911), .B(n4131), .C(n4194), .D(n4195), .Q(n3981) );
  NAND22 U6070 ( .A(n6356), .B(n1449), .Q(n4194) );
  BUF2 U6071 ( .A(n1932), .Q(n6555) );
  BUF2 U6072 ( .A(n1928), .Q(n6573) );
  BUF2 U6073 ( .A(n1926), .Q(n6583) );
  BUF2 U6074 ( .A(n1932), .Q(n6554) );
  BUF2 U6075 ( .A(n1930), .Q(n6563) );
  BUF2 U6076 ( .A(n1926), .Q(n6582) );
  BUF2 U6077 ( .A(n1928), .Q(n6572) );
  BUF2 U6078 ( .A(n1926), .Q(n6581) );
  BUF2 U6079 ( .A(n2015), .Q(n6519) );
  BUF2 U6080 ( .A(n2013), .Q(n6528) );
  BUF2 U6081 ( .A(n2011), .Q(n6536) );
  BUF2 U6082 ( .A(n2015), .Q(n6518) );
  BUF2 U6083 ( .A(n2013), .Q(n6527) );
  BUF2 U6084 ( .A(n2009), .Q(n6545) );
  INV3 U6085 ( .A(n4018), .Q(n1443) );
  INV3 U6086 ( .A(n3368), .Q(n1171) );
  INV3 U6087 ( .A(n3360), .Q(n1174) );
  INV3 U6088 ( .A(n2692), .Q(n1163) );
  INV3 U6089 ( .A(n3361), .Q(n1172) );
  INV3 U6090 ( .A(n2693), .Q(n1165) );
  INV3 U6091 ( .A(n3604), .Q(n1334) );
  BUF2 U6092 ( .A(n1930), .Q(n6564) );
  BUF2 U6093 ( .A(n2011), .Q(n6537) );
  BUF2 U6094 ( .A(n2009), .Q(n6546) );
  INV3 U6095 ( .A(n2700), .Q(n1167) );
  INV3 U6096 ( .A(n6359), .Q(n6360) );
  NOR21 U6097 ( .A(n3361), .B(n6319), .Q(n6359) );
  INV3 U6098 ( .A(n6378), .Q(n6379) );
  NOR21 U6099 ( .A(n3360), .B(n6320), .Q(n6378) );
  NOR21 U6100 ( .A(n2693), .B(n6318), .Q(n2036) );
  BUF2 U6101 ( .A(n3399), .Q(n6358) );
  NOR21 U6102 ( .A(n3365), .B(n6498), .Q(n1943) );
  NOR21 U6103 ( .A(n3364), .B(n6498), .Q(n1944) );
  NOR21 U6104 ( .A(n3365), .B(n6498), .Q(n6404) );
  NOR21 U6105 ( .A(n3364), .B(n6498), .Q(n6409) );
  NOR21 U6106 ( .A(n2697), .B(n6492), .Q(n2026) );
  NOR21 U6107 ( .A(n2696), .B(n6492), .Q(n2027) );
  NOR21 U6108 ( .A(n2697), .B(n6492), .Q(n6468) );
  NOR21 U6109 ( .A(n2696), .B(n6492), .Q(n6473) );
  NOR21 U6110 ( .A(n3364), .B(n6319), .Q(n6385) );
  NOR21 U6111 ( .A(n3364), .B(n6319), .Q(n6384) );
  NOR21 U6112 ( .A(n3364), .B(n6320), .Q(n1945) );
  NOR21 U6113 ( .A(n2696), .B(n6316), .Q(n6448) );
  NOR21 U6114 ( .A(n2696), .B(n6317), .Q(n6447) );
  NOR21 U6115 ( .A(n2696), .B(n6317), .Q(n2028) );
  INV3 U6116 ( .A(n3605), .Q(n1314) );
  BUF2 U6117 ( .A(n1927), .Q(n6577) );
  BUF2 U6118 ( .A(n1925), .Q(n6587) );
  BUF2 U6119 ( .A(n1927), .Q(n6575) );
  BUF2 U6120 ( .A(n1925), .Q(n6585) );
  BUF2 U6121 ( .A(n1927), .Q(n6580) );
  BUF2 U6122 ( .A(n1925), .Q(n6590) );
  BUF2 U6123 ( .A(n1927), .Q(n6579) );
  BUF2 U6124 ( .A(n1925), .Q(n6589) );
  BUF2 U6125 ( .A(n1927), .Q(n6578) );
  BUF2 U6126 ( .A(n1925), .Q(n6588) );
  BUF2 U6127 ( .A(n1927), .Q(n6576) );
  BUF2 U6128 ( .A(n1925), .Q(n6586) );
  BUF2 U6129 ( .A(n1927), .Q(n6574) );
  BUF2 U6130 ( .A(n1925), .Q(n6584) );
  BUF2 U6131 ( .A(n2010), .Q(n6541) );
  BUF2 U6132 ( .A(n2008), .Q(n6550) );
  BUF2 U6133 ( .A(n2010), .Q(n6539) );
  BUF2 U6134 ( .A(n2008), .Q(n6548) );
  BUF2 U6135 ( .A(n2010), .Q(n6544) );
  BUF2 U6136 ( .A(n2008), .Q(n6553) );
  BUF2 U6137 ( .A(n2010), .Q(n6543) );
  BUF2 U6138 ( .A(n2008), .Q(n6552) );
  BUF2 U6139 ( .A(n2010), .Q(n6542) );
  BUF2 U6140 ( .A(n2008), .Q(n6551) );
  BUF2 U6141 ( .A(n2010), .Q(n6540) );
  BUF2 U6142 ( .A(n2008), .Q(n6549) );
  BUF2 U6143 ( .A(n2010), .Q(n6538) );
  BUF2 U6144 ( .A(n2008), .Q(n6547) );
  BUF2 U6145 ( .A(n1931), .Q(n6559) );
  BUF2 U6146 ( .A(n1929), .Q(n6568) );
  BUF2 U6147 ( .A(n1931), .Q(n6557) );
  BUF2 U6148 ( .A(n1929), .Q(n6566) );
  BUF2 U6149 ( .A(n1931), .Q(n6562) );
  BUF2 U6150 ( .A(n1929), .Q(n6571) );
  BUF2 U6151 ( .A(n1931), .Q(n6561) );
  BUF2 U6152 ( .A(n1929), .Q(n6570) );
  BUF2 U6153 ( .A(n1931), .Q(n6560) );
  BUF2 U6154 ( .A(n1929), .Q(n6569) );
  BUF2 U6155 ( .A(n1931), .Q(n6558) );
  BUF2 U6156 ( .A(n1929), .Q(n6567) );
  BUF2 U6157 ( .A(n1931), .Q(n6556) );
  BUF2 U6158 ( .A(n1929), .Q(n6565) );
  BUF2 U6159 ( .A(n2014), .Q(n6523) );
  BUF2 U6160 ( .A(n2012), .Q(n6532) );
  BUF2 U6161 ( .A(n2014), .Q(n6521) );
  BUF2 U6162 ( .A(n2012), .Q(n6530) );
  BUF2 U6163 ( .A(n2014), .Q(n6526) );
  BUF2 U6164 ( .A(n2012), .Q(n6535) );
  BUF2 U6165 ( .A(n2014), .Q(n6525) );
  BUF2 U6166 ( .A(n2012), .Q(n6534) );
  BUF2 U6167 ( .A(n2014), .Q(n6524) );
  BUF2 U6168 ( .A(n2012), .Q(n6533) );
  BUF2 U6169 ( .A(n2014), .Q(n6522) );
  BUF2 U6170 ( .A(n2012), .Q(n6531) );
  BUF2 U6171 ( .A(n2014), .Q(n6520) );
  BUF2 U6172 ( .A(n2012), .Q(n6529) );
  NOR21 U6173 ( .A(n3442), .B(n1363), .Q(n3441) );
  INV3 U6174 ( .A(n3443), .Q(n1363) );
  NOR21 U6175 ( .A(n3360), .B(n6319), .Q(n1952) );
  NOR21 U6176 ( .A(n3368), .B(n6498), .Q(n1954) );
  INV3 U6177 ( .A(n6365), .Q(n6366) );
  NOR21 U6178 ( .A(n3368), .B(n6498), .Q(n6365) );
  INV3 U6179 ( .A(n6422), .Q(n6425) );
  NOR21 U6180 ( .A(n2693), .B(n6316), .Q(n6422) );
  INV3 U6181 ( .A(n6441), .Q(n6444) );
  NOR21 U6182 ( .A(n2692), .B(n6317), .Q(n6441) );
  INV3 U6183 ( .A(n6428), .Q(n6429) );
  NOR21 U6184 ( .A(n2700), .B(n6492), .Q(n6428) );
  NOR21 U6185 ( .A(n2692), .B(n6318), .Q(n6440) );
  NAND22 U6186 ( .A(n1169), .B(n6498), .Q(n1950) );
  NAND22 U6187 ( .A(n1167), .B(n6492), .Q(n2031) );
  INV3 U6188 ( .A(n6394), .Q(n6395) );
  NAND22 U6189 ( .A(n1169), .B(n6498), .Q(n6394) );
  NAND22 U6190 ( .A(n1167), .B(n6492), .Q(n6460) );
  INV3 U6191 ( .A(n6459), .Q(n6461) );
  NAND22 U6192 ( .A(n1167), .B(n6492), .Q(n6459) );
  INV3 U6193 ( .A(n3573), .Q(n1232) );
  NAND31 U6194 ( .A(n1478), .B(n6321), .C(n4064), .Q(n3617) );
  AOI211 U6195 ( .A(n6515), .B(n1411), .C(n6512), .Q(n3658) );
  INV3 U6196 ( .A(n3404), .Q(n6515) );
  AOI211 U6197 ( .A(n6515), .B(n1370), .C(n6512), .Q(n4166) );
  BUF2 U6198 ( .A(n3399), .Q(n6357) );
  AOI211 U6199 ( .A(n3621), .B(n6352), .C(n1413), .Q(n3620) );
  NAND22 U6200 ( .A(n1370), .B(n6210), .Q(n4168) );
  NAND22 U6201 ( .A(n1470), .B(n6348), .Q(n3510) );
  INV3 U6202 ( .A(n1989), .Q(n1494) );
  BUF2 U6203 ( .A(n6593), .Q(n6727) );
  BUF2 U6204 ( .A(n6594), .Q(n6728) );
  BUF2 U6205 ( .A(n6594), .Q(n6729) );
  BUF2 U6206 ( .A(n6595), .Q(n6730) );
  BUF2 U6207 ( .A(n6595), .Q(n6731) );
  BUF2 U6208 ( .A(n6596), .Q(n6732) );
  BUF2 U6209 ( .A(n6596), .Q(n6733) );
  BUF2 U6210 ( .A(n6597), .Q(n6734) );
  BUF2 U6211 ( .A(n6597), .Q(n6735) );
  BUF2 U6212 ( .A(n6598), .Q(n6736) );
  BUF2 U6213 ( .A(n6598), .Q(n6737) );
  BUF2 U6214 ( .A(n6599), .Q(n6738) );
  BUF2 U6215 ( .A(n6599), .Q(n6739) );
  BUF2 U6216 ( .A(n6600), .Q(n6740) );
  BUF2 U6217 ( .A(n6600), .Q(n6741) );
  BUF2 U6218 ( .A(n6601), .Q(n6742) );
  BUF2 U6219 ( .A(n6601), .Q(n6743) );
  BUF2 U6220 ( .A(n6602), .Q(n6744) );
  BUF2 U6221 ( .A(n6602), .Q(n6745) );
  BUF2 U6222 ( .A(n6603), .Q(n6746) );
  BUF2 U6223 ( .A(n6603), .Q(n6747) );
  BUF2 U6224 ( .A(n6604), .Q(n6748) );
  BUF2 U6225 ( .A(n6604), .Q(n6749) );
  BUF2 U6226 ( .A(n6605), .Q(n6750) );
  BUF2 U6227 ( .A(n6605), .Q(n6751) );
  BUF2 U6228 ( .A(n6606), .Q(n6752) );
  BUF2 U6229 ( .A(n6606), .Q(n6753) );
  BUF2 U6230 ( .A(n6607), .Q(n6754) );
  BUF2 U6231 ( .A(n6593), .Q(n6726) );
  BUF2 U6232 ( .A(n6607), .Q(n6755) );
  NOR40 U6233 ( .A(n1364), .B(n3477), .C(n3436), .D(n3467), .Q(n4472) );
  NOR40 U6234 ( .A(n4475), .B(n3907), .C(n3966), .D(n3888), .Q(n4470) );
  NOR40 U6235 ( .A(n4474), .B(n3850), .C(n3832), .D(n3811), .Q(n4471) );
  NOR21 U6236 ( .A(n6269), .B(n1966), .Q(\instruction_decode/reg_MAPP/n1245 )
         );
  NOR21 U6237 ( .A(n6269), .B(n1964), .Q(\instruction_decode/reg_MAPP/n1261 )
         );
  NOR21 U6238 ( .A(n6269), .B(n1965), .Q(\instruction_decode/reg_MAPP/n1253 )
         );
  NOR20 U6239 ( .A(n6269), .B(n1955), .Q(\instruction_decode/reg_MAPP/n1272 )
         );
  NOR21 U6240 ( .A(n1415), .B(n1310), .Q(n4334) );
  NAND22 U6241 ( .A(\instruction_decode/old_ex [3]), .B(n1142), .Q(n1968) );
  NAND22 U6242 ( .A(n6489), .B(\execute/op_21 [23]), .Q(n3843) );
  NOR21 U6243 ( .A(n4542), .B(n4541), .Q(n4404) );
  AOI2111 U6244 ( .A(n1865), .B(n5868), .C(n1981), .D(n1185), .Q(n1978) );
  NOR21 U6245 ( .A(n5945), .B(n5868), .Q(n1981) );
  NAND22 U6246 ( .A(n6489), .B(\execute/op_21 [26]), .Q(n3781) );
  NOR40 U6247 ( .A(n4476), .B(n4176), .C(n4170), .D(n4338), .Q(n4469) );
  NAND31 U6248 ( .A(n1377), .B(n1372), .C(n1374), .Q(n4476) );
  INV3 U6249 ( .A(n4024), .Q(n1381) );
  NOR40 U6250 ( .A(n3398), .B(n3746), .C(n3657), .D(n3718), .Q(n4473) );
  AOI211 U6251 ( .A(n4305), .B(n4306), .C(n4307), .Q(n4303) );
  XNR21 U6252 ( .A(n3735), .B(n3736), .Q(n3734) );
  NAND41 U6253 ( .A(n3709), .B(n3710), .C(n3711), .D(n3712), .Q(
        \execute/old_res [29]) );
  AOI221 U6254 ( .A(n1321), .B(n3720), .C(\execute/alu/sll_175/ML_int[5][29] ), 
        .D(n1353), .Q(n3711) );
  NAND41 U6255 ( .A(n3650), .B(n3651), .C(n3652), .D(n3653), .Q(
        \execute/old_res [30]) );
  AOI211 U6256 ( .A(n1471), .B(n5830), .C(n3674), .Q(n3650) );
  AOI221 U6257 ( .A(n1321), .B(n1292), .C(\execute/alu/sll_175/ML_int[5][30] ), 
        .D(n1353), .Q(n3651) );
  AOI2111 U6258 ( .A(n6513), .B(n3654), .C(n3655), .D(n3656), .Q(n3653) );
  INV3 U6259 ( .A(n4128), .Q(n1372) );
  NAND22 U6260 ( .A(n6489), .B(\execute/op_21 [21]), .Q(n4444) );
  OAI2111 U6261 ( .A(n3407), .B(n3665), .C(n3438), .D(n3666), .Q(n3663) );
  INV3 U6262 ( .A(n3757), .Q(n1408) );
  OAI2111 U6263 ( .A(n4299), .B(n4300), .C(n4301), .D(n4302), .Q(n4298) );
  AOI221 U6264 ( .A(n3721), .B(n6513), .C(n1471), .D(n6346), .Q(n3710) );
  XOR21 U6265 ( .A(n3722), .B(n3723), .Q(n3721) );
  INV3 U6266 ( .A(n3795), .Q(n1404) );
  INV3 U6267 ( .A(n4025), .Q(n1383) );
  INV3 U6268 ( .A(n5829), .Q(n1439) );
  AOI211 U6269 ( .A(n1368), .B(n4318), .C(n4319), .Q(n4317) );
  INV3 U6270 ( .A(n4323), .Q(n1368) );
  INV3 U6271 ( .A(n4111), .Q(n1374) );
  BUF2 U6272 ( .A(n3627), .Q(n6351) );
  INV3 U6273 ( .A(n3777), .Q(n1405) );
  NAND22 U6274 ( .A(n3419), .B(n3398), .Q(n3420) );
  INV3 U6275 ( .A(write_data_reg[0]), .Q(n6931) );
  NAND31 U6276 ( .A(n3727), .B(n3728), .C(n3729), .Q(\execute/old_res [28]) );
  AOI221 U6277 ( .A(\execute/alu/sll_175/ML_int[5][28] ), .B(n1353), .C(n1471), 
        .D(n6345), .Q(n3728) );
  AOI2111 U6278 ( .A(n1457), .B(n3730), .C(n3731), .D(n3732), .Q(n3729) );
  INV3 U6279 ( .A(write_data_reg[4]), .Q(n6940) );
  INV3 U6280 ( .A(n3998), .Q(n1385) );
  INV3 U6281 ( .A(n4083), .Q(n1377) );
  BUF2 U6282 ( .A(n6068), .Q(n6926) );
  INV3 U6283 ( .A(n5830), .Q(n1436) );
  INV3 U6284 ( .A(n4290), .Q(n6338) );
  NOR31 U6285 ( .A(n1491), .B(n1492), .C(n4541), .Q(n4290) );
  INV3 U6286 ( .A(n4542), .Q(n1491) );
  NOR21 U6287 ( .A(n4543), .B(n4541), .Q(n4291) );
  NAND22 U6288 ( .A(n4409), .B(n5946), .Q(n4410) );
  INV3 U6289 ( .A(n3847), .Q(n1392) );
  INV6 U6290 ( .A(n1975), .Q(n1148) );
  NAND22 U6291 ( .A(n6489), .B(\execute/op_21 [30]), .Q(n3659) );
  NOR21 U6292 ( .A(n1963), .B(n1966), .Q(\instruction_decode/reg_MAPP/n1250 )
         );
  NOR21 U6293 ( .A(n1963), .B(n1964), .Q(\instruction_decode/reg_MAPP/n1266 )
         );
  NOR21 U6294 ( .A(n1959), .B(n1966), .Q(\instruction_decode/reg_MAPP/n1246 )
         );
  NOR21 U6295 ( .A(n1957), .B(n1966), .Q(\instruction_decode/reg_MAPP/n1248 )
         );
  NOR21 U6296 ( .A(n1959), .B(n1964), .Q(\instruction_decode/reg_MAPP/n1262 )
         );
  NOR21 U6297 ( .A(n1957), .B(n1964), .Q(\instruction_decode/reg_MAPP/n1264 )
         );
  NOR21 U6298 ( .A(n1959), .B(n1965), .Q(\instruction_decode/reg_MAPP/n1254 )
         );
  NOR21 U6299 ( .A(n1957), .B(n1965), .Q(\instruction_decode/reg_MAPP/n1256 )
         );
  NOR21 U6300 ( .A(n1963), .B(n1965), .Q(\instruction_decode/reg_MAPP/n1258 )
         );
  NAND22 U6301 ( .A(n6489), .B(\execute/op_21 [24]), .Q(n3821) );
  NAND22 U6302 ( .A(n6489), .B(\execute/op_21 [29]), .Q(n3716) );
  NOR21 U6303 ( .A(n1955), .B(n1959), .Q(\instruction_decode/reg_MAPP/n1273 )
         );
  NOR21 U6304 ( .A(n1955), .B(n1957), .Q(\instruction_decode/reg_MAPP/n1275 )
         );
  NOR21 U6305 ( .A(n1955), .B(n1963), .Q(\instruction_decode/reg_MAPP/n1269 )
         );
  NAND22 U6306 ( .A(n6489), .B(\execute/op_21 [25]), .Q(n3793) );
  NAND22 U6307 ( .A(n6489), .B(\execute/op_21 [27]), .Q(n3755) );
  NAND22 U6308 ( .A(n6489), .B(\execute/op_21 [28]), .Q(n3745) );
  NAND41 U6309 ( .A(n3807), .B(n3808), .C(n3809), .D(n3810), .Q(
        \execute/old_res [24]) );
  NAND22 U6310 ( .A(n1452), .B(n3818), .Q(n3808) );
  NAND41 U6311 ( .A(n3748), .B(n3749), .C(n3750), .D(n3751), .Q(
        \execute/old_res [27]) );
  AOI221 U6312 ( .A(\execute/alu/sll_175/ML_int[5][27] ), .B(n1353), .C(n6236), 
        .D(n1240), .Q(n3750) );
  NAND41 U6313 ( .A(n3787), .B(n3788), .C(n3789), .D(n3790), .Q(
        \execute/old_res [25]) );
  AOI221 U6314 ( .A(n1321), .B(n3797), .C(\execute/alu/sll_175/ML_int[5][25] ), 
        .D(n1353), .Q(n3789) );
  NAND41 U6315 ( .A(n3675), .B(n3676), .C(n3677), .D(n3678), .Q(
        \execute/old_res [2]) );
  NAND22 U6316 ( .A(n1349), .B(n3705), .Q(n3676) );
  NAND41 U6317 ( .A(n3882), .B(n3883), .C(n3884), .D(n3885), .Q(
        \execute/old_res [21]) );
  AOI221 U6318 ( .A(n3859), .B(n3546), .C(\execute/alu/sll_175/ML_int[5][21] ), 
        .D(n1353), .Q(n3884) );
  NAND41 U6319 ( .A(n3828), .B(n3829), .C(n3830), .D(n3831), .Q(
        \execute/old_res [23]) );
  NAND22 U6320 ( .A(n1451), .B(n3839), .Q(n3829) );
  NAND41 U6321 ( .A(n3767), .B(n3768), .C(n3769), .D(n3770), .Q(
        \execute/old_res [26]) );
  AOI2111 U6322 ( .A(n1471), .B(n1428), .C(n3771), .D(n3772), .Q(n3770) );
  NAND41 U6323 ( .A(n3900), .B(n3901), .C(n3902), .D(n3903), .Q(
        \execute/old_res [20]) );
  NAND22 U6324 ( .A(n3919), .B(n6515), .Q(n3901) );
  XNR21 U6325 ( .A(n3844), .B(n3845), .Q(n3841) );
  XNR21 U6326 ( .A(n3823), .B(n3824), .Q(n3822) );
  AOI221 U6327 ( .A(n3783), .B(n1470), .C(n6513), .D(n3784), .Q(n3767) );
  AOI221 U6328 ( .A(n3859), .B(n3519), .C(n6236), .D(n3498), .Q(n3858) );
  XNR21 U6329 ( .A(n3868), .B(n3869), .Q(n3857) );
  AOI2111 U6330 ( .A(n1448), .B(n3904), .C(n3905), .D(n3906), .Q(n3903) );
  AOI221 U6331 ( .A(n3760), .B(n6513), .C(n1471), .D(n6344), .Q(n3749) );
  XNR21 U6332 ( .A(n3761), .B(n3762), .Q(n3760) );
  BUF2 U6333 ( .A(n1468), .Q(n6323) );
  INV3 U6334 ( .A(n6980), .Q(n6979) );
  BUF2 U6335 ( .A(n1468), .Q(n6324) );
  INV3 U6336 ( .A(write_data_reg[1]), .Q(n6933) );
  INV3 U6337 ( .A(write_data_reg[2]), .Q(n6935) );
  BUF2 U6338 ( .A(n6929), .Q(n6927) );
  INV3 U6339 ( .A(n4413), .Q(n1481) );
  NOR21 U6340 ( .A(n4163), .B(n4164), .Q(n4162) );
  BUF2 U6341 ( .A(n6929), .Q(n6928) );
  NAND22 U6342 ( .A(n3388), .B(n1247), .Q(\execute/old_res [9]) );
  INV3 U6343 ( .A(n3389), .Q(n1247) );
  AOI2111 U6344 ( .A(n6512), .B(n3398), .C(n3405), .D(n3406), .Q(n3388) );
  OAI2111 U6345 ( .A(n3390), .B(n3391), .C(n3392), .D(n3393), .Q(n3389) );
  INV3 U6346 ( .A(n1866), .Q(n1141) );
  NAND22 U6347 ( .A(n6489), .B(\execute/op_21 [31]), .Q(n3622) );
  NOR21 U6348 ( .A(n1961), .B(n1966), .Q(\instruction_decode/reg_MAPP/n1252 )
         );
  NOR21 U6349 ( .A(n1961), .B(n1964), .Q(\instruction_decode/reg_MAPP/n1268 )
         );
  NOR21 U6350 ( .A(n1961), .B(n1965), .Q(\instruction_decode/reg_MAPP/n1260 )
         );
  NOR21 U6351 ( .A(n1955), .B(n1961), .Q(\instruction_decode/reg_MAPP/n1271 )
         );
  NOR21 U6352 ( .A(n1955), .B(n1958), .Q(\instruction_decode/reg_MAPP/n1274 )
         );
  NOR21 U6353 ( .A(n1955), .B(n1956), .Q(\instruction_decode/reg_MAPP/n1276 )
         );
  NOR21 U6354 ( .A(n1955), .B(n1962), .Q(\instruction_decode/reg_MAPP/n1270 )
         );
  NOR21 U6355 ( .A(n1958), .B(n1965), .Q(\instruction_decode/reg_MAPP/n1255 )
         );
  NOR21 U6356 ( .A(n1962), .B(n1965), .Q(\instruction_decode/reg_MAPP/n1259 )
         );
  NOR21 U6357 ( .A(n1956), .B(n1965), .Q(\instruction_decode/reg_MAPP/n1257 )
         );
  NOR21 U6358 ( .A(n1962), .B(n1964), .Q(\instruction_decode/reg_MAPP/n1267 )
         );
  NOR21 U6359 ( .A(n1956), .B(n1964), .Q(\instruction_decode/reg_MAPP/n1265 )
         );
  NOR21 U6360 ( .A(n1958), .B(n1964), .Q(\instruction_decode/reg_MAPP/n1263 )
         );
  NOR21 U6361 ( .A(n1962), .B(n1966), .Q(\instruction_decode/reg_MAPP/n1251 )
         );
  NOR21 U6362 ( .A(n1956), .B(n1966), .Q(\instruction_decode/reg_MAPP/n1249 )
         );
  NOR21 U6363 ( .A(n1958), .B(n1966), .Q(\instruction_decode/reg_MAPP/n1247 )
         );
  NOR40 U6364 ( .A(n4485), .B(n1393), .C(n1370), .D(n1367), .Q(n4484) );
  AOI2111 U6365 ( .A(n3527), .B(n6513), .C(n3556), .D(n6512), .Q(n3555) );
  NAND22 U6366 ( .A(n1476), .B(n4282), .Q(n4395) );
  XNR21 U6367 ( .A(n3996), .B(n3997), .Q(n3988) );
  NOR40 U6368 ( .A(n4513), .B(n1358), .C(n1401), .D(n1398), .Q(n4482) );
  NAND41 U6369 ( .A(n3456), .B(n3457), .C(n3458), .D(n3459), .Q(
        \execute/old_res [7]) );
  OAI311 U6370 ( .A(n3478), .B(n3479), .C(n1276), .D(n1473), .Q(n3457) );
  NAND41 U6371 ( .A(n4179), .B(n4180), .C(n4181), .D(n4182), .Q(
        \execute/old_res [11]) );
  AOI2111 U6372 ( .A(n1321), .B(n3481), .C(n4203), .D(n4204), .Q(n4181) );
  NOR40 U6373 ( .A(n4183), .B(n4184), .C(n4185), .D(n4186), .Q(n4182) );
  NAND41 U6374 ( .A(n3488), .B(n3489), .C(n3490), .D(n1236), .Q(
        \execute/old_res [6]) );
  NAND22 U6375 ( .A(n4207), .B(n4208), .Q(n3484) );
  NAND22 U6376 ( .A(n4211), .B(n4212), .Q(n3481) );
  NOR40 U6377 ( .A(n4526), .B(n1410), .C(n1409), .D(n1411), .Q(n4481) );
  NAND22 U6378 ( .A(n4266), .B(n4267), .Q(n3518) );
  NAND22 U6379 ( .A(n4268), .B(n4269), .Q(n3499) );
  XNR21 U6380 ( .A(n4214), .B(n4215), .Q(n4213) );
  AOI2111 U6381 ( .A(n1336), .B(n3469), .C(n3597), .D(n3598), .Q(n3595) );
  NAND31 U6382 ( .A(n3959), .B(n3960), .C(n3961), .Q(\execute/old_res [19]) );
  AOI2111 U6383 ( .A(n1447), .B(n3962), .C(n3963), .D(n3964), .Q(n3961) );
  NAND31 U6384 ( .A(n3424), .B(n3425), .C(n3426), .Q(\execute/old_res [8]) );
  NAND22 U6385 ( .A(n4346), .B(n4347), .Q(n3574) );
  NAND22 U6386 ( .A(n4396), .B(n4397), .Q(n3571) );
  NAND22 U6387 ( .A(n4348), .B(n4349), .Q(n4178) );
  NAND22 U6388 ( .A(n4144), .B(n4145), .Q(n3545) );
  AOI211 U6389 ( .A(n3396), .B(n1313), .C(n3397), .Q(n3392) );
  OAI311 U6390 ( .A(n3398), .B(n1427), .C(n6357), .D(n3400), .Q(n3397) );
  NAND22 U6391 ( .A(n1427), .B(n1365), .Q(n3400) );
  INV3 U6392 ( .A(n3401), .Q(n1365) );
  NAND22 U6393 ( .A(n3955), .B(n3956), .Q(n3536) );
  INV3 U6394 ( .A(n6992), .Q(n6991) );
  INV3 U6395 ( .A(n6986), .Q(n6985) );
  INV3 U6396 ( .A(n6968), .Q(n6967) );
  INV3 U6397 ( .A(n6990), .Q(n6989) );
  INV3 U6398 ( .A(n6988), .Q(n6987) );
  INV3 U6399 ( .A(n6982), .Q(n6981) );
  INV3 U6400 ( .A(n6950), .Q(n6949) );
  INV3 U6401 ( .A(n4281), .Q(n1476) );
  INV3 U6402 ( .A(n4408), .Q(n1493) );
  NAND22 U6403 ( .A(n3547), .B(n3548), .Q(\execute/old_res [4]) );
  NOR40 U6404 ( .A(n3549), .B(n3550), .C(n3551), .D(n3552), .Q(n3548) );
  NOR40 U6405 ( .A(n3565), .B(n3566), .C(n3567), .D(n3568), .Q(n3547) );
  NAND31 U6406 ( .A(n4366), .B(n3564), .C(n4367), .Q(n3390) );
  NAND22 U6407 ( .A(n4281), .B(n4282), .Q(n3407) );
  INV3 U6408 ( .A(n3693), .Q(n1309) );
  NAND22 U6409 ( .A(n3357), .B(n3358), .Q(n1932) );
  NAND22 U6410 ( .A(n4142), .B(n4143), .Q(n3394) );
  INV3 U6411 ( .A(n4189), .Q(n1244) );
  NAND22 U6412 ( .A(n4190), .B(n4191), .Q(n4189) );
  NAND22 U6413 ( .A(n4205), .B(n4206), .Q(n3460) );
  NAND22 U6414 ( .A(n4373), .B(n4374), .Q(n3427) );
  NAND22 U6415 ( .A(n4252), .B(n4253), .Q(n3502) );
  INV3 U6416 ( .A(n4375), .Q(n1233) );
  NAND22 U6417 ( .A(n4376), .B(n4377), .Q(n4375) );
  INV3 U6418 ( .A(n3469), .Q(n1253) );
  NAND22 U6419 ( .A(n4257), .B(n4258), .Q(n3500) );
  AOI2111 U6420 ( .A(n1314), .B(n3573), .C(n4368), .D(n4369), .Q(n4365) );
  NAND22 U6421 ( .A(n3946), .B(n3947), .Q(n3423) );
  NOR21 U6422 ( .A(n1849), .B(n6089), .Q(n1851) );
  BUF2 U6423 ( .A(\instruction_decode/hazard_unit/n5 ), .Q(n6762) );
  INV3 U6424 ( .A(n3943), .Q(n1252) );
  NAND22 U6425 ( .A(n2689), .B(n2688), .Q(n2010) );
  NAND22 U6426 ( .A(n2686), .B(n2688), .Q(n2008) );
  NAND22 U6427 ( .A(n3357), .B(n3356), .Q(n1927) );
  NAND22 U6428 ( .A(n3354), .B(n3356), .Q(n1925) );
  NAND22 U6429 ( .A(n2689), .B(n2691), .Q(n2014) );
  NAND22 U6430 ( .A(n2686), .B(n2691), .Q(n2012) );
  NAND22 U6431 ( .A(n3357), .B(n3359), .Q(n1931) );
  NAND22 U6432 ( .A(n3354), .B(n3359), .Q(n1929) );
  NAND22 U6433 ( .A(n2704), .B(n2688), .Q(n2696) );
  NAND22 U6434 ( .A(n3372), .B(n3356), .Q(n3364) );
  NAND22 U6435 ( .A(n3359), .B(n3370), .Q(n3361) );
  NAND22 U6436 ( .A(n3356), .B(n3370), .Q(n3368) );
  NAND22 U6437 ( .A(n3358), .B(n3370), .Q(n3360) );
  NAND22 U6438 ( .A(n2691), .B(n2702), .Q(n2693) );
  NAND22 U6439 ( .A(n2688), .B(n2702), .Q(n2700) );
  NAND22 U6440 ( .A(n2690), .B(n2702), .Q(n2692) );
  NAND22 U6441 ( .A(n3357), .B(n3355), .Q(n1928) );
  NAND22 U6442 ( .A(n3354), .B(n3355), .Q(n1926) );
  NAND22 U6443 ( .A(n2689), .B(n2687), .Q(n2011) );
  NAND22 U6444 ( .A(n2686), .B(n2687), .Q(n2009) );
  NAND22 U6445 ( .A(n3354), .B(n3358), .Q(n1930) );
  NAND22 U6446 ( .A(n2689), .B(n2690), .Q(n2015) );
  NAND22 U6447 ( .A(n2686), .B(n2690), .Q(n2013) );
  NAND22 U6448 ( .A(n3355), .B(n3370), .Q(n3365) );
  NAND22 U6449 ( .A(n2687), .B(n2702), .Q(n2697) );
  NOR21 U6450 ( .A(inst_out[24]), .B(inst_out[22]), .Q(n3372) );
  NOR21 U6451 ( .A(inst_out[18]), .B(inst_out[16]), .Q(n2691) );
  NOR21 U6452 ( .A(inst_out[23]), .B(inst_out[21]), .Q(n3359) );
  NOR21 U6453 ( .A(inst_out[19]), .B(inst_out[17]), .Q(n2704) );
  NAND22 U6454 ( .A(n4378), .B(n4379), .Q(n3573) );
  INV3 U6455 ( .A(n3371), .Q(n1169) );
  NAND22 U6456 ( .A(n3372), .B(n3355), .Q(n3371) );
  INV3 U6457 ( .A(n2703), .Q(n1161) );
  NAND22 U6458 ( .A(n2704), .B(n2687), .Q(n2703) );
  INV3 U6459 ( .A(n3373), .Q(n1175) );
  NAND22 U6460 ( .A(n3358), .B(n3372), .Q(n3373) );
  INV3 U6461 ( .A(n2705), .Q(n1164) );
  NAND22 U6462 ( .A(n2690), .B(n2704), .Q(n2705) );
  AOI2111 U6463 ( .A(n3402), .B(n3398), .C(n3403), .D(n6512), .Q(n3401) );
  NOR21 U6464 ( .A(n3398), .B(n6514), .Q(n3403) );
  INV3 U6465 ( .A(n4343), .Q(n1478) );
  BUF2 U6466 ( .A(n6501), .Q(n6499) );
  BUF2 U6467 ( .A(inst_out[25]), .Q(n6500) );
  BUF2 U6468 ( .A(n6495), .Q(n6493) );
  BUF2 U6469 ( .A(inst_out[20]), .Q(n6494) );
  INV3 U6470 ( .A(n6346), .Q(n1434) );
  BUF2 U6471 ( .A(inst_out[25]), .Q(n6501) );
  BUF2 U6472 ( .A(inst_out[20]), .Q(n6495) );
  NAND22 U6473 ( .A(n5945), .B(n6085), .Q(n1972) );
  INV3 U6474 ( .A(n1771), .Q(n1185) );
  INV3 U6475 ( .A(n1980), .Q(n1187) );
  INV3 U6476 ( .A(n1854), .Q(n1465) );
  BUF2 U6477 ( .A(n1108), .Q(n6594) );
  BUF2 U6478 ( .A(n1108), .Q(n6595) );
  BUF2 U6479 ( .A(n1108), .Q(n6596) );
  BUF2 U6480 ( .A(n1108), .Q(n6597) );
  BUF2 U6481 ( .A(n1108), .Q(n6598) );
  BUF2 U6482 ( .A(n1108), .Q(n6599) );
  BUF2 U6483 ( .A(n1108), .Q(n6600) );
  BUF2 U6484 ( .A(n1108), .Q(n6601) );
  BUF2 U6485 ( .A(n1108), .Q(n6602) );
  BUF2 U6486 ( .A(n1108), .Q(n6603) );
  BUF2 U6487 ( .A(n1108), .Q(n6604) );
  BUF2 U6488 ( .A(n1108), .Q(n6605) );
  BUF2 U6489 ( .A(n1108), .Q(n6606) );
  BUF2 U6490 ( .A(n1108), .Q(n6607) );
  BUF2 U6491 ( .A(n1108), .Q(n6593) );
  NOR21 U6492 ( .A(n6246), .B(n6247), .Q(n4419) );
  NAND22 U6493 ( .A(n4509), .B(n4510), .Q(n3998) );
  AOI221 U6494 ( .A(ram_adr[18]), .B(n6336), .C(n6339), .D(data_1[18]), .Q(
        n4510) );
  AOI221 U6495 ( .A(n6503), .B(write_data_reg[18]), .C(pc_ex[18]), .D(n6324), 
        .Q(n4509) );
  NAND22 U6496 ( .A(n4531), .B(n4532), .Q(n3718) );
  AOI221 U6497 ( .A(ram_adr[29]), .B(n6336), .C(n6339), .D(data_1[29]), .Q(
        n4532) );
  AOI221 U6498 ( .A(n6503), .B(write_data_reg[29]), .C(pc_ex[29]), .D(n6324), 
        .Q(n4531) );
  NAND22 U6499 ( .A(n4514), .B(n4515), .Q(n3832) );
  AOI221 U6500 ( .A(ram_adr[23]), .B(n6336), .C(n6339), .D(data_1[23]), .Q(
        n4515) );
  AOI221 U6501 ( .A(n6503), .B(write_data_reg[23]), .C(pc_ex[23]), .D(n6324), 
        .Q(n4514) );
  NAND22 U6502 ( .A(n4518), .B(n4519), .Q(n3477) );
  NAND22 U6503 ( .A(n4535), .B(n4536), .Q(n3467) );
  AOI221 U6504 ( .A(ram_adr[7]), .B(n6336), .C(n6339), .D(data_1[7]), .Q(n4536) );
  AOI221 U6505 ( .A(n6503), .B(n6945), .C(pc_ex[7]), .D(n6324), .Q(n4535) );
  NAND22 U6506 ( .A(n4516), .B(n4517), .Q(n3811) );
  XNR21 U6507 ( .A(write_register_ex[2]), .B(rs[2]), .Q(n4553) );
  XNR21 U6508 ( .A(write_register_ex[0]), .B(rs[0]), .Q(n4552) );
  NOR31 U6509 ( .A(n4555), .B(n4556), .C(n4557), .Q(n4554) );
  XNR21 U6510 ( .A(pc_rom[30]), .B(n1851), .Q(n1850) );
  NAND22 U6511 ( .A(n4494), .B(n4495), .Q(n4083) );
  AOI221 U6512 ( .A(n6504), .B(n6961), .C(pc_ex[15]), .D(n6323), .Q(n4494) );
  AOI221 U6513 ( .A(ram_adr[15]), .B(n6337), .C(n6340), .D(data_1[15]), .Q(
        n4495) );
  NAND22 U6514 ( .A(n1851), .B(pc_rom[30]), .Q(n1864) );
  NAND22 U6515 ( .A(n4501), .B(n4502), .Q(n3966) );
  AOI221 U6516 ( .A(n6504), .B(write_data_reg[19]), .C(pc_ex[19]), .D(n6324), 
        .Q(n4501) );
  AOI221 U6517 ( .A(ram_adr[19]), .B(n6336), .C(n6340), .D(data_1[19]), .Q(
        n4502) );
  NAND22 U6518 ( .A(n4490), .B(n4491), .Q(n3907) );
  AOI221 U6519 ( .A(n6504), .B(write_data_reg[20]), .C(pc_ex[20]), .D(n6323), 
        .Q(n4490) );
  AOI221 U6520 ( .A(ram_adr[20]), .B(n6337), .C(n6340), .D(data_1[20]), .Q(
        n4491) );
  NAND22 U6521 ( .A(n4507), .B(n4508), .Q(n3777) );
  NAND22 U6522 ( .A(n4527), .B(n4528), .Q(n3657) );
  NAND22 U6523 ( .A(n4492), .B(n4493), .Q(n4111) );
  NAND22 U6524 ( .A(n4522), .B(n4523), .Q(n3757) );
  NAND22 U6525 ( .A(n4524), .B(n4525), .Q(n3795) );
  NAND22 U6526 ( .A(n4503), .B(n4504), .Q(n3888) );
  INV3 U6527 ( .A(write_data_reg[3]), .Q(n6938) );
  NAND22 U6528 ( .A(n4529), .B(n4530), .Q(n3746) );
  NAND31 U6529 ( .A(n5848), .B(n5941), .C(n5867), .Q(n1960) );
  NAND22 U6530 ( .A(n4498), .B(n4499), .Q(n4176) );
  NAND22 U6531 ( .A(n4402), .B(n4403), .Q(n3542) );
  INV3 U6532 ( .A(inst_rom[2]), .Q(n1138) );
  AOI221 U6533 ( .A(n6437), .B(n5913), .C(n6440), .D(n6046), .Q(n2186) );
  AOI221 U6534 ( .A(n6426), .B(n6026), .C(n5534), .D(n6432), .Q(n2185) );
  AOI221 U6535 ( .A(n6374), .B(n5931), .C(n6383), .D(n6060), .Q(n3169) );
  AOI2111 U6536 ( .A(n6391), .B(n5428), .C(n3187), .D(n3188), .Q(n3170) );
  AOI221 U6537 ( .A(n6437), .B(n6021), .C(n6445), .D(n5932), .Q(n2165) );
  AOI221 U6538 ( .A(n2036), .B(n6022), .C(n5542), .D(n6432), .Q(n2164) );
  AOI2111 U6539 ( .A(n5544), .B(n6452), .C(n2183), .D(n2184), .Q(n2166) );
  AOI221 U6540 ( .A(n6437), .B(n5911), .C(n6440), .D(n6044), .Q(n2228) );
  AOI221 U6541 ( .A(n2036), .B(n6024), .C(n5518), .D(n6432), .Q(n2227) );
  AOI2111 U6542 ( .A(n5520), .B(n6450), .C(n2246), .D(n2247), .Q(n2229) );
  AOI221 U6543 ( .A(n6438), .B(n5912), .C(n6445), .D(n6045), .Q(n2249) );
  AOI221 U6544 ( .A(n2036), .B(n6025), .C(n5510), .D(n6433), .Q(n2248) );
  AOI2111 U6545 ( .A(n5512), .B(n6449), .C(n2267), .D(n2268), .Q(n2250) );
  AOI221 U6546 ( .A(n2034), .B(n5914), .C(n6443), .D(n6047), .Q(n2270) );
  AOI221 U6547 ( .A(n6423), .B(n6027), .C(n5502), .D(n6431), .Q(n2269) );
  AOI2111 U6548 ( .A(n5504), .B(n6452), .C(n2288), .D(n2289), .Q(n2271) );
  AOI221 U6549 ( .A(n6438), .B(n5909), .C(n6442), .D(n6042), .Q(n2291) );
  AOI221 U6550 ( .A(n2036), .B(n5908), .C(n5494), .D(n6431), .Q(n2290) );
  AOI2111 U6551 ( .A(n5496), .B(n6451), .C(n2309), .D(n2310), .Q(n2292) );
  AOI221 U6552 ( .A(n6436), .B(n5915), .C(n6443), .D(n6048), .Q(n2312) );
  AOI221 U6553 ( .A(n6424), .B(n6028), .C(n5486), .D(n6430), .Q(n2311) );
  AOI2111 U6554 ( .A(n5488), .B(n6454), .C(n2330), .D(n2331), .Q(n2313) );
  AOI221 U6555 ( .A(n6436), .B(n5861), .C(n6442), .D(n5937), .Q(n2333) );
  AOI221 U6556 ( .A(n6423), .B(n5862), .C(n5478), .D(n6431), .Q(n2332) );
  AOI2111 U6557 ( .A(n5480), .B(n6453), .C(n2351), .D(n2352), .Q(n2334) );
  AOI221 U6558 ( .A(n6436), .B(n6030), .C(n6442), .D(n5933), .Q(n2459) );
  AOI221 U6559 ( .A(n6423), .B(n6031), .C(n5434), .D(n6430), .Q(n2458) );
  AOI2111 U6560 ( .A(n5436), .B(n6449), .C(n2477), .D(n2478), .Q(n2460) );
  AOI221 U6561 ( .A(n6436), .B(n5859), .C(n6446), .D(n5934), .Q(n2501) );
  AOI221 U6562 ( .A(n6423), .B(n6032), .C(n5418), .D(n6431), .Q(n2500) );
  AOI2111 U6563 ( .A(n5420), .B(n6453), .C(n2519), .D(n2520), .Q(n2502) );
  AOI221 U6564 ( .A(n6439), .B(n5917), .C(n6445), .D(n6049), .Q(n2522) );
  AOI221 U6565 ( .A(n6426), .B(n5918), .C(n5410), .D(n6433), .Q(n2521) );
  AOI2111 U6566 ( .A(n5412), .B(n6450), .C(n2540), .D(n2541), .Q(n2523) );
  AOI221 U6567 ( .A(n6438), .B(n5919), .C(n6445), .D(n6050), .Q(n2543) );
  AOI221 U6568 ( .A(n2036), .B(n5920), .C(n5402), .D(n6433), .Q(n2542) );
  AOI2111 U6569 ( .A(n5404), .B(n6449), .C(n2561), .D(n2562), .Q(n2544) );
  AOI221 U6570 ( .A(n6437), .B(n5921), .C(n6440), .D(n6051), .Q(n2564) );
  AOI221 U6571 ( .A(n2036), .B(n6033), .C(n5394), .D(n6432), .Q(n2563) );
  AOI2111 U6572 ( .A(n5396), .B(n6452), .C(n2582), .D(n2583), .Q(n2565) );
  AOI221 U6573 ( .A(n2034), .B(n5922), .C(n6443), .D(n6052), .Q(n2606) );
  AOI221 U6574 ( .A(n6423), .B(n6034), .C(n5378), .D(n6431), .Q(n2605) );
  AOI2111 U6575 ( .A(n5380), .B(n6450), .C(n2624), .D(n2625), .Q(n2607) );
  AOI221 U6576 ( .A(n6439), .B(n5923), .C(n6442), .D(n6053), .Q(n2627) );
  AOI221 U6577 ( .A(n6424), .B(n5924), .C(n5370), .D(n6431), .Q(n2626) );
  AOI2111 U6578 ( .A(n5372), .B(n6449), .C(n2645), .D(n2646), .Q(n2628) );
  AOI221 U6579 ( .A(n6436), .B(n5925), .C(n6443), .D(n6054), .Q(n2648) );
  AOI221 U6580 ( .A(n6424), .B(n6035), .C(n5362), .D(n6430), .Q(n2647) );
  AOI2111 U6581 ( .A(n5364), .B(n6449), .C(n2666), .D(n2667), .Q(n2649) );
  AOI221 U6582 ( .A(n6438), .B(n5926), .C(n6446), .D(n6056), .Q(n2102) );
  AOI221 U6583 ( .A(n6426), .B(n5927), .C(n5566), .D(n6433), .Q(n2101) );
  AOI2111 U6584 ( .A(n5568), .B(n6454), .C(n2120), .D(n2121), .Q(n2103) );
  AOI221 U6585 ( .A(n6438), .B(n5928), .C(n6445), .D(n6057), .Q(n2123) );
  AOI221 U6586 ( .A(n2036), .B(n6036), .C(n5558), .D(n6433), .Q(n2122) );
  AOI2111 U6587 ( .A(n5560), .B(n6453), .C(n2141), .D(n2142), .Q(n2124) );
  AOI221 U6588 ( .A(n6437), .B(n5929), .C(n6442), .D(n6058), .Q(n2144) );
  AOI221 U6589 ( .A(n2036), .B(n6037), .C(n5550), .D(n6432), .Q(n2143) );
  AOI2111 U6590 ( .A(n5552), .B(n6453), .C(n2162), .D(n2163), .Q(n2145) );
  AOI221 U6591 ( .A(n6438), .B(n5910), .C(n6440), .D(n6043), .Q(n2207) );
  AOI221 U6592 ( .A(n2036), .B(n6023), .C(n5526), .D(n6433), .Q(n2206) );
  AOI2111 U6593 ( .A(n5528), .B(n6451), .C(n2225), .D(n2226), .Q(n2208) );
  AOI221 U6594 ( .A(n2034), .B(n5930), .C(n6443), .D(n6059), .Q(n2438) );
  AOI221 U6595 ( .A(n6424), .B(n6038), .C(n5442), .D(n6431), .Q(n2437) );
  AOI2111 U6596 ( .A(n5352), .B(n6450), .C(n2456), .D(n2457), .Q(n2439) );
  AOI221 U6597 ( .A(n6436), .B(n5843), .C(n6443), .D(n5935), .Q(n2669) );
  AOI221 U6598 ( .A(n6423), .B(n6039), .C(n5358), .D(n6430), .Q(n2668) );
  AOI2111 U6599 ( .A(n6454), .B(n6020), .C(n2698), .D(n2699), .Q(n2670) );
  AOI221 U6600 ( .A(n6372), .B(n5844), .C(n6383), .D(n5936), .Q(n1912) );
  AOI221 U6601 ( .A(n6364), .B(n5860), .C(n5386), .D(n6370), .Q(n1911) );
  AOI2111 U6602 ( .A(n5388), .B(n6389), .C(n1946), .D(n1947), .Q(n1913) );
  AOI221 U6603 ( .A(n6439), .B(n5863), .C(n6446), .D(n5938), .Q(n2354) );
  AOI221 U6604 ( .A(n6427), .B(n6040), .C(n5470), .D(n6433), .Q(n2353) );
  AOI2111 U6605 ( .A(n5472), .B(n6452), .C(n2372), .D(n2373), .Q(n2355) );
  AOI221 U6606 ( .A(n2034), .B(n5834), .C(n6440), .D(n6061), .Q(n2375) );
  AOI221 U6607 ( .A(n2036), .B(n5836), .C(n5462), .D(n6432), .Q(n2374) );
  AOI2111 U6608 ( .A(n5464), .B(n6451), .C(n2393), .D(n2394), .Q(n2376) );
  AOI221 U6609 ( .A(n6439), .B(n5837), .C(n6442), .D(n5850), .Q(n2396) );
  AOI221 U6610 ( .A(n6427), .B(n5864), .C(n5454), .D(n6430), .Q(n2395) );
  AOI2111 U6611 ( .A(n5456), .B(n6451), .C(n2414), .D(n2415), .Q(n2397) );
  AOI221 U6612 ( .A(n6439), .B(n6029), .C(n6446), .D(n5849), .Q(n2417) );
  AOI221 U6613 ( .A(n6427), .B(n5916), .C(n5446), .D(n6430), .Q(n2416) );
  AOI2111 U6614 ( .A(n5448), .B(n6450), .C(n2435), .D(n2436), .Q(n2418) );
  AOI221 U6615 ( .A(n6439), .B(n5845), .C(n6446), .D(n5865), .Q(n1995) );
  AOI221 U6616 ( .A(n6427), .B(n6041), .C(n5598), .D(n6430), .Q(n1994) );
  AOI2111 U6617 ( .A(n5600), .B(n6454), .C(n2029), .D(n2030), .Q(n1996) );
  AOI221 U6618 ( .A(n6436), .B(n5833), .C(n6445), .D(n5835), .Q(n2039) );
  AOI221 U6619 ( .A(n6424), .B(n5838), .C(n5590), .D(n6431), .Q(n2038) );
  AOI2111 U6620 ( .A(n5592), .B(n6453), .C(n2057), .D(n2058), .Q(n2040) );
  AOI221 U6621 ( .A(n6439), .B(n5846), .C(n6446), .D(n5866), .Q(n2060) );
  AOI221 U6622 ( .A(n6423), .B(n5847), .C(n5582), .D(n6430), .Q(n2059) );
  AOI2111 U6623 ( .A(n5584), .B(n6450), .C(n2078), .D(n2079), .Q(n2061) );
  AOI221 U6624 ( .A(n6439), .B(n5841), .C(n6446), .D(n6055), .Q(n2081) );
  AOI221 U6625 ( .A(n6427), .B(n5842), .C(n5574), .D(n6430), .Q(n2080) );
  AOI2111 U6626 ( .A(n5576), .B(n6449), .C(n2099), .D(n2100), .Q(n2082) );
  AOI221 U6627 ( .A(n6372), .B(n5909), .C(n6380), .D(n6042), .Q(n2980) );
  AOI221 U6628 ( .A(n6376), .B(n6021), .C(n6381), .D(n5932), .Q(n2854) );
  AOI221 U6629 ( .A(n6362), .B(n6022), .C(n5542), .D(n6369), .Q(n2853) );
  AOI221 U6630 ( .A(n6376), .B(n5910), .C(n6381), .D(n6043), .Q(n2896) );
  AOI221 U6631 ( .A(n6362), .B(n6023), .C(n5526), .D(n1954), .Q(n2895) );
  AOI221 U6632 ( .A(n6372), .B(n5911), .C(n1952), .D(n6044), .Q(n2917) );
  AOI221 U6633 ( .A(n6361), .B(n6024), .C(n5518), .D(n6369), .Q(n2916) );
  AOI221 U6634 ( .A(n6375), .B(n5912), .C(n6380), .D(n6045), .Q(n2938) );
  AOI221 U6635 ( .A(n6361), .B(n6025), .C(n5510), .D(n6367), .Q(n2937) );
  AOI221 U6636 ( .A(n6376), .B(n5913), .C(n6382), .D(n6046), .Q(n2875) );
  AOI221 U6637 ( .A(n6362), .B(n6026), .C(n5534), .D(n1954), .Q(n2874) );
  AOI221 U6638 ( .A(n6372), .B(n5914), .C(n6383), .D(n6047), .Q(n2959) );
  AOI221 U6639 ( .A(n6363), .B(n6027), .C(n5502), .D(n6370), .Q(n2958) );
  AOI2111 U6640 ( .A(n5504), .B(n6390), .C(n2977), .D(n2978), .Q(n2960) );
  AOI221 U6641 ( .A(n6374), .B(n5915), .C(n6380), .D(n6048), .Q(n3001) );
  AOI221 U6642 ( .A(n6361), .B(n6028), .C(n5486), .D(n6368), .Q(n3000) );
  AOI2111 U6643 ( .A(n5488), .B(n6390), .C(n3019), .D(n3020), .Q(n3002) );
  AOI221 U6644 ( .A(n6375), .B(n6029), .C(n6380), .D(n5849), .Q(n3106) );
  AOI221 U6645 ( .A(n6363), .B(n5916), .C(n5446), .D(n6368), .Q(n3105) );
  AOI2111 U6646 ( .A(n5448), .B(n6387), .C(n3124), .D(n3125), .Q(n3107) );
  AOI221 U6647 ( .A(n6377), .B(n6030), .C(n6383), .D(n5933), .Q(n3148) );
  AOI221 U6648 ( .A(n6364), .B(n6031), .C(n5434), .D(n6367), .Q(n3147) );
  AOI2111 U6649 ( .A(n5436), .B(n6391), .C(n3166), .D(n3167), .Q(n3149) );
  AOI221 U6650 ( .A(n6376), .B(n5859), .C(n6382), .D(n5934), .Q(n3190) );
  AOI221 U6651 ( .A(n6362), .B(n6032), .C(n5418), .D(n6370), .Q(n3189) );
  AOI2111 U6652 ( .A(n5420), .B(n6390), .C(n3208), .D(n3209), .Q(n3191) );
  AOI221 U6653 ( .A(n6372), .B(n5917), .C(n6382), .D(n6049), .Q(n3211) );
  AOI221 U6654 ( .A(n6361), .B(n5918), .C(n5410), .D(n6369), .Q(n3210) );
  AOI2111 U6655 ( .A(n5412), .B(n6387), .C(n3229), .D(n3230), .Q(n3212) );
  AOI221 U6656 ( .A(n6377), .B(n5919), .C(n6381), .D(n6050), .Q(n3232) );
  AOI221 U6657 ( .A(n6363), .B(n5920), .C(n5402), .D(n1954), .Q(n3231) );
  AOI2111 U6658 ( .A(n5404), .B(n6386), .C(n3250), .D(n3251), .Q(n3233) );
  AOI221 U6659 ( .A(n6377), .B(n5921), .C(n1952), .D(n6051), .Q(n3253) );
  AOI221 U6660 ( .A(n6361), .B(n6033), .C(n5394), .D(n6369), .Q(n3252) );
  AOI2111 U6661 ( .A(n5396), .B(n6389), .C(n3271), .D(n3272), .Q(n3254) );
  AOI221 U6662 ( .A(n6375), .B(n5922), .C(n6380), .D(n6052), .Q(n3274) );
  AOI221 U6663 ( .A(n6363), .B(n6034), .C(n5378), .D(n6368), .Q(n3273) );
  AOI2111 U6664 ( .A(n5380), .B(n6388), .C(n3292), .D(n3293), .Q(n3275) );
  AOI221 U6665 ( .A(n6372), .B(n5923), .C(n6383), .D(n6053), .Q(n3295) );
  AOI221 U6666 ( .A(n6363), .B(n5924), .C(n5370), .D(n6368), .Q(n3294) );
  AOI2111 U6667 ( .A(n5372), .B(n6387), .C(n3313), .D(n3314), .Q(n3296) );
  AOI221 U6668 ( .A(n6372), .B(n5925), .C(n6383), .D(n6054), .Q(n3316) );
  AOI221 U6669 ( .A(n6363), .B(n6035), .C(n5362), .D(n6367), .Q(n3315) );
  AOI2111 U6670 ( .A(n5364), .B(n6386), .C(n3334), .D(n3335), .Q(n3317) );
  AOI221 U6671 ( .A(n6376), .B(n5841), .C(n6381), .D(n6055), .Q(n2770) );
  AOI221 U6672 ( .A(n6362), .B(n5842), .C(n5574), .D(n6369), .Q(n2769) );
  AOI2111 U6673 ( .A(n5576), .B(n6391), .C(n2788), .D(n2789), .Q(n2771) );
  AOI221 U6674 ( .A(n6372), .B(n5926), .C(n6382), .D(n6056), .Q(n2791) );
  AOI221 U6675 ( .A(n6361), .B(n5927), .C(n5566), .D(n6368), .Q(n2790) );
  AOI2111 U6676 ( .A(n5568), .B(n6390), .C(n2809), .D(n2810), .Q(n2792) );
  AOI221 U6677 ( .A(n6377), .B(n5928), .C(n6381), .D(n6057), .Q(n2812) );
  AOI221 U6678 ( .A(n6361), .B(n6036), .C(n5558), .D(n6370), .Q(n2811) );
  AOI2111 U6679 ( .A(n5560), .B(n6387), .C(n2830), .D(n2831), .Q(n2813) );
  AOI221 U6680 ( .A(n6377), .B(n5929), .C(n1952), .D(n6058), .Q(n2833) );
  AOI221 U6681 ( .A(n6361), .B(n6037), .C(n5550), .D(n6367), .Q(n2832) );
  AOI2111 U6682 ( .A(n5552), .B(n6386), .C(n2851), .D(n2852), .Q(n2834) );
  AOI221 U6683 ( .A(n6372), .B(n5930), .C(n6380), .D(n6059), .Q(n3127) );
  AOI221 U6684 ( .A(n6364), .B(n6038), .C(n5442), .D(n6367), .Q(n3126) );
  AOI2111 U6685 ( .A(n5352), .B(n6386), .C(n3145), .D(n3146), .Q(n3128) );
  AOI221 U6686 ( .A(n6374), .B(n5843), .C(n6383), .D(n5935), .Q(n3337) );
  AOI221 U6687 ( .A(n6363), .B(n6039), .C(n5358), .D(n6368), .Q(n3336) );
  AOI2111 U6688 ( .A(n6390), .B(n6020), .C(n3366), .D(n3367), .Q(n3338) );
  AOI221 U6689 ( .A(n6436), .B(n5931), .C(n6443), .D(n6060), .Q(n2480) );
  AOI221 U6690 ( .A(n6424), .B(n5940), .C(n5426), .D(n6430), .Q(n2479) );
  AOI2111 U6691 ( .A(n5428), .B(n6454), .C(n2498), .D(n2499), .Q(n2481) );
  AOI221 U6692 ( .A(n6436), .B(n5844), .C(n6445), .D(n5936), .Q(n2585) );
  AOI221 U6693 ( .A(n2036), .B(n5860), .C(n5386), .D(n6433), .Q(n2584) );
  AOI2111 U6694 ( .A(n5388), .B(n6451), .C(n2603), .D(n2604), .Q(n2586) );
  AOI221 U6695 ( .A(n6372), .B(n5861), .C(n6383), .D(n5937), .Q(n3022) );
  AOI221 U6696 ( .A(n6364), .B(n5862), .C(n5478), .D(n6370), .Q(n3021) );
  AOI2111 U6697 ( .A(n5480), .B(n6389), .C(n3040), .D(n3041), .Q(n3023) );
  AOI221 U6698 ( .A(n6377), .B(n5863), .C(n6383), .D(n5938), .Q(n3043) );
  AOI221 U6699 ( .A(n6363), .B(n6040), .C(n5470), .D(n6370), .Q(n3042) );
  AOI2111 U6700 ( .A(n5472), .B(n6388), .C(n3061), .D(n3062), .Q(n3044) );
  AOI221 U6701 ( .A(n6372), .B(n5834), .C(n6383), .D(n6061), .Q(n3064) );
  AOI221 U6702 ( .A(n6364), .B(n5836), .C(n5462), .D(n6368), .Q(n3063) );
  AOI2111 U6703 ( .A(n5464), .B(n6389), .C(n3082), .D(n3083), .Q(n3065) );
  AOI221 U6704 ( .A(n6372), .B(n5837), .C(n6383), .D(n5850), .Q(n3085) );
  AOI221 U6705 ( .A(n6364), .B(n5864), .C(n5454), .D(n6370), .Q(n3084) );
  AOI2111 U6706 ( .A(n5456), .B(n6388), .C(n3103), .D(n3104), .Q(n3086) );
  AOI221 U6707 ( .A(n6377), .B(n5845), .C(n6383), .D(n5865), .Q(n2707) );
  AOI221 U6708 ( .A(n6363), .B(n6041), .C(n5598), .D(n6367), .Q(n2706) );
  AOI2111 U6709 ( .A(n5600), .B(n6388), .C(n2725), .D(n2726), .Q(n2708) );
  AOI221 U6710 ( .A(n6377), .B(n5833), .C(n1952), .D(n5835), .Q(n2728) );
  AOI221 U6711 ( .A(n6363), .B(n5838), .C(n5590), .D(n6369), .Q(n2727) );
  AOI2111 U6712 ( .A(n5592), .B(n6387), .C(n2746), .D(n2747), .Q(n2729) );
  AOI221 U6713 ( .A(n6377), .B(n5846), .C(n6383), .D(n5866), .Q(n2749) );
  AOI221 U6714 ( .A(n6363), .B(n5847), .C(n5582), .D(n1954), .Q(n2748) );
  AOI2111 U6715 ( .A(n5584), .B(n6386), .C(n2767), .D(n2768), .Q(n2750) );
  NAND22 U6716 ( .A(n4486), .B(n4487), .Q(n4170) );
  AOI221 U6717 ( .A(n6504), .B(n6953), .C(pc_ex[11]), .D(n6323), .Q(n4486) );
  AOI221 U6718 ( .A(ram_adr[11]), .B(n6337), .C(n6340), .D(data_1[11]), .Q(
        n4487) );
  NOR21 U6719 ( .A(n1255), .B(n5611), .Q(n5767) );
  NOR21 U6720 ( .A(n1255), .B(n5608), .Q(n5768) );
  NAND22 U6721 ( .A(n4520), .B(n4521), .Q(n3850) );
  AOI221 U6722 ( .A(n6503), .B(n6975), .C(pc_ex[22]), .D(n6323), .Q(n4520) );
  AOI221 U6723 ( .A(ram_adr[22]), .B(n6337), .C(n6339), .D(data_1[22]), .Q(
        n4521) );
  OAI311 U6724 ( .A(n5868), .B(n5715), .C(n5718), .D(n6085), .Q(n1984) );
  NAND31 U6725 ( .A(n5696), .B(n5697), .C(n5695), .Q(n1992) );
  NAND22 U6726 ( .A(n4537), .B(n4538), .Q(n3436) );
  AOI221 U6727 ( .A(n6503), .B(n6947), .C(pc_ex[8]), .D(n6324), .Q(n4537) );
  AOI221 U6728 ( .A(ram_adr[8]), .B(n6337), .C(n6339), .D(data_1[8]), .Q(n4538) );
  NAND22 U6729 ( .A(n4511), .B(n4512), .Q(n4025) );
  NOR40 U6730 ( .A(n3161), .B(n3162), .C(n3163), .D(n3164), .Q(n3155) );
  NOR40 U6731 ( .A(n3245), .B(n3246), .C(n3247), .D(n3248), .Q(n3239) );
  NOR40 U6732 ( .A(n2367), .B(n2368), .C(n2369), .D(n2370), .Q(n2361) );
  NOR40 U6733 ( .A(n2409), .B(n2410), .C(n2411), .D(n2412), .Q(n2403) );
  NOR40 U6734 ( .A(n2430), .B(n2431), .C(n2432), .D(n2433), .Q(n2424) );
  NOR40 U6735 ( .A(n2472), .B(n2473), .C(n2474), .D(n2475), .Q(n2466) );
  NOR40 U6736 ( .A(n2535), .B(n2536), .C(n2537), .D(n2538), .Q(n2529) );
  NOR40 U6737 ( .A(n2556), .B(n2557), .C(n2558), .D(n2559), .Q(n2550) );
  NOR40 U6738 ( .A(n2577), .B(n2578), .C(n2579), .D(n2580), .Q(n2571) );
  NOR40 U6739 ( .A(n2640), .B(n2641), .C(n2642), .D(n2643), .Q(n2634) );
  NOR40 U6740 ( .A(n2661), .B(n2662), .C(n2663), .D(n2664), .Q(n2655) );
  NOR40 U6741 ( .A(n2052), .B(n2053), .C(n2054), .D(n2055), .Q(n2046) );
  NOR40 U6742 ( .A(n2073), .B(n2074), .C(n2075), .D(n2076), .Q(n2067) );
  AOI221 U6743 ( .A(n6332), .B(data_2[4]), .C(n5816), .D(ram_adr[4]), .Q(n4433) );
  NOR21 U6744 ( .A(n5604), .B(n1255), .Q(n5772) );
  NOR21 U6745 ( .A(n5605), .B(n1255), .Q(n5771) );
  NOR21 U6746 ( .A(n5606), .B(n1255), .Q(n5770) );
  NOR21 U6747 ( .A(n5607), .B(n1255), .Q(n5769) );
  AOI211 U6748 ( .A(n5716), .B(n1865), .C(n1185), .Q(n1982) );
  XNR21 U6749 ( .A(n6067), .B(write_register[1]), .Q(n4565) );
  NOR41 U6750 ( .A(n1492), .B(n5823), .C(n4550), .D(n4551), .Q(n4548) );
  NOR40 U6751 ( .A(n2525), .B(n2526), .C(n2527), .D(n2528), .Q(n2524) );
  NOR40 U6752 ( .A(n2609), .B(n2610), .C(n2611), .D(n2612), .Q(n2608) );
  NOR40 U6753 ( .A(n3235), .B(n3236), .C(n3237), .D(n3238), .Q(n3234) );
  NOR40 U6754 ( .A(n3298), .B(n3299), .C(n3300), .D(n3301), .Q(n3297) );
  NOR40 U6755 ( .A(n2630), .B(n2631), .C(n2632), .D(n2633), .Q(n2629) );
  INV3 U6756 ( .A(\instruction_decode/N13 ), .Q(n1158) );
  XNR21 U6757 ( .A(n1799), .B(pc_rom[5]), .Q(n1798) );
  XNR21 U6758 ( .A(n1831), .B(pc_rom[27]), .Q(n1830) );
  XNR21 U6759 ( .A(n1828), .B(pc_rom[25]), .Q(n1827) );
  XNR21 U6760 ( .A(n1790), .B(pc_rom[17]), .Q(n1789) );
  XOR31 U6761 ( .A(n6263), .B(inst_out[13]), .C(
        \instruction_decode/add_358/carry [15]), .Q(n6262) );
  NAND22 U6762 ( .A(n4488), .B(n4489), .Q(n4338) );
  INV3 U6763 ( .A(\instruction_decode/N15 ), .Q(n1157) );
  XNR21 U6764 ( .A(n1862), .B(pc_rom[7]), .Q(n1861) );
  XOR21 U6765 ( .A(rs[1]), .B(write_register_ex[1]), .Q(n4557) );
  XNR21 U6766 ( .A(n6089), .B(n1849), .Q(n1848) );
  NAND22 U6767 ( .A(n4496), .B(n4497), .Q(n4128) );
  INV3 U6768 ( .A(inst_rom[20]), .Q(n1120) );
  BUF6 U6769 ( .A(n3939), .Q(n6341) );
  OAI2111 U6770 ( .A(n6931), .B(n6505), .C(n4477), .D(n4478), .Q(n3939) );
  AOI221 U6771 ( .A(n1467), .B(n5944), .C(pc_ex[0]), .D(n6324), .Q(n4478) );
  AOI221 U6772 ( .A(ram_adr[0]), .B(n6336), .C(n6340), .D(data_1[0]), .Q(n4477) );
  NAND22 U6773 ( .A(n4505), .B(n4506), .Q(n4024) );
  XNR21 U6774 ( .A(n1793), .B(pc_rom[23]), .Q(n1792) );
  XNR21 U6775 ( .A(n1825), .B(pc_rom[21]), .Q(n1824) );
  XNR21 U6776 ( .A(n1787), .B(pc_rom[19]), .Q(n1786) );
  INV3 U6777 ( .A(\instruction_decode/N21 ), .Q(n1154) );
  INV3 U6778 ( .A(\instruction_decode/N19 ), .Q(n1155) );
  XNR21 U6779 ( .A(n1834), .B(pc_rom[11]), .Q(n1833) );
  INV3 U6780 ( .A(\instruction_decode/N17 ), .Q(n1156) );
  XNR21 U6781 ( .A(n1796), .B(pc_rom[9]), .Q(n1795) );
  INV3 U6782 ( .A(\instruction_decode/N12 ), .Q(n1159) );
  XOR21 U6783 ( .A(pc_rom[4]), .B(n1784), .Q(n1783) );
  XNR21 U6784 ( .A(n4581), .B(n5701), .Q(n1812) );
  AOI221 U6785 ( .A(n1142), .B(inst_out[1]), .C(\instruction_decode/N11 ), .D(
        n1143), .Q(n1813) );
  XNR21 U6786 ( .A(pc_rom[20]), .B(n1844), .Q(n1842) );
  AOI221 U6787 ( .A(n1142), .B(inst_out[18]), .C(pc_out[20]), .D(n1143), .Q(
        n1843) );
  XNR21 U6788 ( .A(pc_rom[22]), .B(n1808), .Q(n1806) );
  AOI221 U6789 ( .A(n1142), .B(n6491), .C(pc_out[22]), .D(n1143), .Q(n1807) );
  XNR21 U6790 ( .A(pc_rom[16]), .B(n1805), .Q(n1803) );
  AOI221 U6791 ( .A(n1142), .B(inst_out[14]), .C(pc_out[16]), .D(n1143), .Q(
        n1804) );
  XNR21 U6792 ( .A(pc_rom[14]), .B(n1822), .Q(n1820) );
  AOI221 U6793 ( .A(n1142), .B(inst_out[12]), .C(\instruction_decode/N22 ), 
        .D(n1143), .Q(n1821) );
  XNR21 U6794 ( .A(pc_rom[12]), .B(n1819), .Q(n1817) );
  AOI221 U6795 ( .A(n1142), .B(inst_out[10]), .C(\instruction_decode/N20 ), 
        .D(n1143), .Q(n1818) );
  XNR21 U6796 ( .A(pc_rom[10]), .B(n1837), .Q(n1835) );
  AOI221 U6797 ( .A(n1142), .B(inst_out[8]), .C(\instruction_decode/N18 ), .D(
        n1143), .Q(n1836) );
  XNR21 U6798 ( .A(pc_rom[8]), .B(n1859), .Q(n1857) );
  AOI221 U6799 ( .A(n1142), .B(inst_out[6]), .C(\instruction_decode/N16 ), .D(
        n1143), .Q(n1858) );
  XNR21 U6800 ( .A(pc_rom[6]), .B(n1802), .Q(n1800) );
  AOI221 U6801 ( .A(n1142), .B(inst_out[4]), .C(\instruction_decode/N14 ), .D(
        n1143), .Q(n1801) );
  XNR21 U6802 ( .A(pc_rom[24]), .B(n1847), .Q(n1845) );
  AOI221 U6803 ( .A(n1142), .B(inst_out[22]), .C(pc_out[24]), .D(n1143), .Q(
        n1846) );
  XNR21 U6804 ( .A(pc_rom[26]), .B(n1811), .Q(n1809) );
  AOI221 U6805 ( .A(n1142), .B(inst_out[24]), .C(pc_out[26]), .D(n1143), .Q(
        n1810) );
  XNR21 U6806 ( .A(pc_rom[18]), .B(n1776), .Q(n1774) );
  AOI221 U6807 ( .A(n1142), .B(inst_out[16]), .C(pc_out[18]), .D(n1143), .Q(
        n1775) );
  AOI221 U6808 ( .A(n5543), .B(n6406), .C(n5540), .D(n6411), .Q(n2871) );
  AOI221 U6809 ( .A(n5535), .B(n6405), .C(n5532), .D(n6410), .Q(n2892) );
  AOI221 U6810 ( .A(n5519), .B(n6405), .C(n5516), .D(n6410), .Q(n2934) );
  AOI221 U6811 ( .A(n5511), .B(n6407), .C(n5508), .D(n6412), .Q(n2955) );
  AOI221 U6812 ( .A(n5503), .B(n6406), .C(n5500), .D(n6411), .Q(n2976) );
  AOI221 U6813 ( .A(n5495), .B(n6405), .C(n5492), .D(n6410), .Q(n2997) );
  AOI221 U6814 ( .A(n5471), .B(n6407), .C(n5468), .D(n6412), .Q(n3060) );
  AOI221 U6815 ( .A(n5463), .B(n6406), .C(n5460), .D(n6411), .Q(n3081) );
  AOI221 U6816 ( .A(n5455), .B(n6407), .C(n5452), .D(n6412), .Q(n3102) );
  AOI221 U6817 ( .A(n5447), .B(n6405), .C(n5444), .D(n6410), .Q(n3123) );
  AOI221 U6818 ( .A(n5435), .B(n6407), .C(n5432), .D(n6412), .Q(n3165) );
  AOI221 U6819 ( .A(n5419), .B(n6406), .C(n5416), .D(n6411), .Q(n3207) );
  AOI221 U6820 ( .A(n5411), .B(n6406), .C(n5408), .D(n6411), .Q(n3228) );
  AOI221 U6821 ( .A(n5403), .B(n6405), .C(n5400), .D(n6410), .Q(n3249) );
  AOI221 U6822 ( .A(n5379), .B(n6405), .C(n5376), .D(n6410), .Q(n3291) );
  AOI221 U6823 ( .A(n5371), .B(n6407), .C(n5368), .D(n6412), .Q(n3312) );
  AOI221 U6824 ( .A(n5363), .B(n6406), .C(n5360), .D(n6411), .Q(n3333) );
  AOI221 U6825 ( .A(n5599), .B(n6407), .C(n5596), .D(n6412), .Q(n2724) );
  AOI221 U6826 ( .A(n5591), .B(n6406), .C(n5588), .D(n6411), .Q(n2745) );
  AOI221 U6827 ( .A(n5583), .B(n6407), .C(n5580), .D(n6412), .Q(n2766) );
  AOI221 U6828 ( .A(n5575), .B(n6405), .C(n5572), .D(n6410), .Q(n2787) );
  AOI221 U6829 ( .A(n5559), .B(n6407), .C(n5556), .D(n6412), .Q(n2829) );
  AOI221 U6830 ( .A(n5551), .B(n6406), .C(n5548), .D(n6411), .Q(n2850) );
  AOI221 U6831 ( .A(n5359), .B(n6405), .C(n5356), .D(n6410), .Q(n3363) );
  AOI221 U6832 ( .A(n5543), .B(n6469), .C(n5540), .D(n6474), .Q(n2182) );
  AOI221 U6833 ( .A(n5535), .B(n6472), .C(n5532), .D(n6477), .Q(n2203) );
  AOI221 U6834 ( .A(n5519), .B(n6470), .C(n5516), .D(n6475), .Q(n2245) );
  AOI221 U6835 ( .A(n5511), .B(n6469), .C(n5508), .D(n6474), .Q(n2266) );
  AOI221 U6836 ( .A(n5503), .B(n6472), .C(n5500), .D(n6477), .Q(n2287) );
  AOI221 U6837 ( .A(n5495), .B(n6471), .C(n5492), .D(n6476), .Q(n2308) );
  AOI221 U6838 ( .A(n5487), .B(n6470), .C(n5484), .D(n6475), .Q(n2329) );
  AOI221 U6839 ( .A(n5479), .B(n6469), .C(n5476), .D(n6474), .Q(n2350) );
  AOI221 U6840 ( .A(n5471), .B(n6472), .C(n5468), .D(n6477), .Q(n2371) );
  AOI221 U6841 ( .A(n5463), .B(n6471), .C(n5460), .D(n6476), .Q(n2392) );
  AOI221 U6842 ( .A(n5455), .B(n6470), .C(n5452), .D(n6475), .Q(n2413) );
  AOI221 U6843 ( .A(n5447), .B(n6469), .C(n5444), .D(n6474), .Q(n2434) );
  AOI221 U6844 ( .A(n5435), .B(n6471), .C(n5432), .D(n6476), .Q(n2476) );
  AOI221 U6845 ( .A(n5427), .B(n6470), .C(n5424), .D(n6475), .Q(n2497) );
  AOI221 U6846 ( .A(n5419), .B(n6469), .C(n5416), .D(n6474), .Q(n2518) );
  AOI221 U6847 ( .A(n5411), .B(n6472), .C(n5408), .D(n6477), .Q(n2539) );
  AOI221 U6848 ( .A(n5403), .B(n6471), .C(n5400), .D(n6476), .Q(n2560) );
  AOI221 U6849 ( .A(n5395), .B(n6470), .C(n5392), .D(n6475), .Q(n2581) );
  AOI221 U6850 ( .A(n5387), .B(n6469), .C(n5384), .D(n6474), .Q(n2602) );
  AOI221 U6851 ( .A(n5379), .B(n6472), .C(n5376), .D(n6477), .Q(n2623) );
  AOI221 U6852 ( .A(n5363), .B(n6470), .C(n5360), .D(n6475), .Q(n2665) );
  AOI221 U6853 ( .A(n5599), .B(n6472), .C(n5596), .D(n6477), .Q(n2025) );
  AOI221 U6854 ( .A(n5591), .B(n6471), .C(n5588), .D(n6476), .Q(n2056) );
  AOI221 U6855 ( .A(n5583), .B(n6470), .C(n5580), .D(n6475), .Q(n2077) );
  AOI221 U6856 ( .A(n5575), .B(n6469), .C(n5572), .D(n6474), .Q(n2098) );
  AOI221 U6857 ( .A(n5567), .B(n6472), .C(n5564), .D(n6477), .Q(n2119) );
  AOI221 U6858 ( .A(n5559), .B(n6471), .C(n5556), .D(n6476), .Q(n2140) );
  AOI221 U6859 ( .A(n5551), .B(n6470), .C(n5548), .D(n6475), .Q(n2161) );
  AOI221 U6860 ( .A(n5527), .B(n6471), .C(n5524), .D(n6476), .Q(n2224) );
  AOI221 U6861 ( .A(n5443), .B(n6472), .C(n5440), .D(n6477), .Q(n2455) );
  AOI221 U6862 ( .A(n5359), .B(n6469), .C(n5356), .D(n6474), .Q(n2695) );
  AOI221 U6863 ( .A(n5487), .B(n6408), .C(n5484), .D(n6413), .Q(n3018) );
  AOI221 U6864 ( .A(n5479), .B(n6408), .C(n5476), .D(n6413), .Q(n3039) );
  AOI221 U6865 ( .A(n5395), .B(n6408), .C(n5392), .D(n6413), .Q(n3270) );
  AOI221 U6866 ( .A(n5387), .B(n6408), .C(n5384), .D(n6413), .Q(n1942) );
  AOI221 U6867 ( .A(n5567), .B(n6408), .C(n5564), .D(n6413), .Q(n2808) );
  AOI221 U6868 ( .A(n5527), .B(n6408), .C(n5524), .D(n6413), .Q(n2913) );
  AOI221 U6869 ( .A(n5443), .B(n6408), .C(n5440), .D(n6413), .Q(n3144) );
  NOR31 U6870 ( .A(n6216), .B(n5700), .C(n1992), .Q(n4544) );
  NOR21 U6871 ( .A(n6282), .B(n1139), .Q(n5765) );
  INV3 U6872 ( .A(inst_rom[1]), .Q(n1139) );
  NOR21 U6873 ( .A(n6285), .B(n1128), .Q(n5754) );
  INV3 U6874 ( .A(inst_rom[12]), .Q(n1128) );
  NOR21 U6875 ( .A(n6282), .B(n1129), .Q(n5755) );
  INV3 U6876 ( .A(inst_rom[11]), .Q(n1129) );
  INV3 U6877 ( .A(inst_rom[3]), .Q(n1137) );
  INV3 U6878 ( .A(inst_rom[23]), .Q(n1117) );
  INV3 U6879 ( .A(inst_rom[15]), .Q(n1125) );
  NOR21 U6880 ( .A(n6293), .B(n1124), .Q(n5750) );
  INV3 U6881 ( .A(inst_rom[16]), .Q(n1124) );
  NOR21 U6882 ( .A(n6291), .B(n1126), .Q(n5752) );
  INV3 U6883 ( .A(inst_rom[14]), .Q(n1126) );
  NOR21 U6884 ( .A(n6301), .B(n1127), .Q(n5753) );
  INV3 U6885 ( .A(inst_rom[13]), .Q(n1127) );
  NAND22 U6886 ( .A(n5710), .B(n1968), .Q(\instruction_decode/old_rd [4]) );
  NAND22 U6887 ( .A(n5711), .B(n1968), .Q(\instruction_decode/old_rd [3]) );
  NAND22 U6888 ( .A(n5714), .B(n1968), .Q(\instruction_decode/old_rd [2]) );
  NAND22 U6889 ( .A(n5712), .B(n1968), .Q(\instruction_decode/old_rd [1]) );
  NAND22 U6890 ( .A(n5713), .B(n1968), .Q(\instruction_decode/old_rd [0]) );
  NOR21 U6891 ( .A(n6302), .B(n1112), .Q(n5738) );
  INV3 U6892 ( .A(inst_rom[28]), .Q(n1112) );
  NOR21 U6893 ( .A(n6303), .B(n1135), .Q(n5761) );
  INV3 U6894 ( .A(inst_rom[5]), .Q(n1135) );
  NOR21 U6895 ( .A(n6303), .B(n1136), .Q(n5762) );
  INV3 U6896 ( .A(inst_rom[4]), .Q(n1136) );
  NOR21 U6897 ( .A(n6302), .B(n1121), .Q(n5747) );
  INV3 U6898 ( .A(inst_rom[19]), .Q(n1121) );
  NOR21 U6899 ( .A(n6294), .B(n1130), .Q(n5756) );
  INV3 U6900 ( .A(inst_rom[10]), .Q(n1130) );
  NOR21 U6901 ( .A(n6291), .B(n1131), .Q(n5757) );
  INV3 U6902 ( .A(inst_rom[9]), .Q(n1131) );
  NOR21 U6903 ( .A(n6306), .B(n1132), .Q(n5758) );
  INV3 U6904 ( .A(inst_rom[8]), .Q(n1132) );
  NOR21 U6905 ( .A(n6294), .B(n1111), .Q(n5737) );
  INV3 U6906 ( .A(inst_rom[29]), .Q(n1111) );
  NOR21 U6907 ( .A(n6306), .B(n1133), .Q(n5759) );
  INV3 U6908 ( .A(inst_rom[7]), .Q(n1133) );
  NOR21 U6909 ( .A(n6305), .B(n1134), .Q(n5760) );
  INV3 U6910 ( .A(inst_rom[6]), .Q(n1134) );
  NOR21 U6911 ( .A(n6305), .B(n1109), .Q(n5735) );
  INV3 U6912 ( .A(inst_rom[31]), .Q(n1109) );
  NOR21 U6913 ( .A(n6293), .B(n1110), .Q(n5736) );
  INV3 U6914 ( .A(inst_rom[30]), .Q(n1110) );
  NOR21 U6915 ( .A(n6291), .B(n1116), .Q(n5742) );
  INV3 U6916 ( .A(inst_rom[24]), .Q(n1116) );
  NOR21 U6917 ( .A(n6288), .B(n1119), .Q(n5745) );
  INV3 U6918 ( .A(inst_rom[21]), .Q(n1119) );
  NOR21 U6919 ( .A(n6292), .B(n1114), .Q(n5740) );
  INV3 U6920 ( .A(inst_rom[26]), .Q(n1114) );
  NOR21 U6921 ( .A(n6293), .B(n1113), .Q(n5739) );
  INV3 U6922 ( .A(inst_rom[27]), .Q(n1113) );
  NOR21 U6923 ( .A(n6293), .B(n1118), .Q(n5744) );
  INV3 U6924 ( .A(inst_rom[22]), .Q(n1118) );
  NOR21 U6925 ( .A(n6301), .B(n1122), .Q(n5748) );
  INV3 U6926 ( .A(inst_rom[18]), .Q(n1122) );
  NOR21 U6927 ( .A(n6294), .B(n1123), .Q(n5749) );
  INV3 U6928 ( .A(inst_rom[17]), .Q(n1123) );
  NOR21 U6929 ( .A(n6301), .B(n1140), .Q(n5766) );
  INV3 U6930 ( .A(inst_rom[0]), .Q(n1140) );
  NOR21 U6931 ( .A(n6291), .B(n1115), .Q(n5741) );
  INV3 U6932 ( .A(inst_rom[25]), .Q(n1115) );
  AOI211 U6933 ( .A(n6085), .B(n1185), .C(n1977), .Q(n1976) );
  AOI211 U6934 ( .A(n1972), .B(n1771), .C(n5716), .Q(n1977) );
  INV3 U6935 ( .A(write_data_reg[11]), .Q(n6954) );
  INV3 U6936 ( .A(write_data_reg[5]), .Q(n6942) );
  NAND22 U6937 ( .A(n4539), .B(n4540), .Q(n1991) );
  NAND31 U6938 ( .A(n5715), .B(n6085), .C(n6279), .Q(n1969) );
  AOI211 U6939 ( .A(n1769), .B(n1151), .C(n6085), .Q(n5773) );
  INV3 U6940 ( .A(n1770), .Q(n1151) );
  AOI221 U6941 ( .A(n5371), .B(n6471), .C(n5368), .D(n6476), .Q(n2644) );
  INV3 U6942 ( .A(write_data_reg[22]), .Q(n6976) );
  INV3 U6943 ( .A(write_data_reg[21]), .Q(n6974) );
  INV3 U6944 ( .A(write_data_reg[20]), .Q(n6972) );
  INV3 U6945 ( .A(write_data_reg[19]), .Q(n6970) );
  INV3 U6946 ( .A(write_data_reg[17]), .Q(n6966) );
  INV3 U6947 ( .A(write_data_reg[16]), .Q(n6964) );
  INV3 U6948 ( .A(write_data_reg[15]), .Q(n6962) );
  INV3 U6949 ( .A(write_data_reg[12]), .Q(n6956) );
  INV3 U6950 ( .A(write_data_reg[7]), .Q(n6946) );
  INV3 U6951 ( .A(write_data_reg[6]), .Q(n6944) );
  INV3 U6952 ( .A(write_data_reg[10]), .Q(n6952) );
  INV3 U6953 ( .A(write_data_reg[13]), .Q(n6958) );
  INV3 U6954 ( .A(write_data_reg[24]), .Q(n6980) );
  INV3 U6955 ( .A(write_data_reg[23]), .Q(n6978) );
  INV3 U6956 ( .A(write_data_reg[26]), .Q(n6984) );
  INV3 U6957 ( .A(write_data_reg[8]), .Q(n6948) );
  INV3 U6958 ( .A(write_data_reg[14]), .Q(n6960) );
  INV3 U6959 ( .A(write_data_reg[31]), .Q(n6994) );
  NOR40 U6960 ( .A(n3382), .B(n3383), .C(n3384), .D(n3385), .Q(n3374) );
  NOR40 U6961 ( .A(n3376), .B(n3377), .C(n3378), .D(n3379), .Q(n3375) );
  NOR21 U6962 ( .A(inst_out[23]), .B(n5725), .Q(n3358) );
  NOR21 U6963 ( .A(inst_out[22]), .B(n5721), .Q(n3357) );
  NAND22 U6964 ( .A(n1811), .B(pc_rom[26]), .Q(n1831) );
  NAND22 U6965 ( .A(n1776), .B(pc_rom[18]), .Q(n1787) );
  NAND22 U6966 ( .A(pc_rom[22]), .B(n1808), .Q(n1793) );
  NAND22 U6967 ( .A(pc_rom[28]), .B(n1853), .Q(n1849) );
  NAND22 U6968 ( .A(pc_rom[20]), .B(n1844), .Q(n1825) );
  NAND22 U6969 ( .A(pc_rom[24]), .B(n1847), .Q(n1828) );
  NAND22 U6970 ( .A(pc_rom[4]), .B(n1784), .Q(n1799) );
  NAND22 U6971 ( .A(pc_rom[12]), .B(n1819), .Q(n1781) );
  NAND22 U6972 ( .A(pc_rom[14]), .B(n1822), .Q(n1816) );
  NAND22 U6973 ( .A(pc_rom[16]), .B(n1805), .Q(n1790) );
  NAND22 U6974 ( .A(pc_rom[10]), .B(n1837), .Q(n1834) );
  NAND22 U6975 ( .A(pc_rom[8]), .B(n1859), .Q(n1796) );
  NAND22 U6976 ( .A(pc_rom[6]), .B(n1802), .Q(n1862) );
  NOR21 U6977 ( .A(n4581), .B(n5701), .Q(n1784) );
  NOR21 U6978 ( .A(n6076), .B(n1834), .Q(n1819) );
  NOR21 U6979 ( .A(n6078), .B(n1781), .Q(n1822) );
  NOR21 U6980 ( .A(n6079), .B(n1816), .Q(n1805) );
  NOR21 U6981 ( .A(n6077), .B(n1796), .Q(n1837) );
  NOR21 U6982 ( .A(n6070), .B(n1862), .Q(n1859) );
  NOR21 U6983 ( .A(n6083), .B(n1825), .Q(n1808) );
  NOR21 U6984 ( .A(n6071), .B(n1799), .Q(n1802) );
  NOR21 U6985 ( .A(n1793), .B(n6087), .Q(n1847) );
  NOR21 U6986 ( .A(n1787), .B(n6082), .Q(n1844) );
  NOR21 U6987 ( .A(n5729), .B(n6080), .Q(\instruction_decode/add_358/carry [3]) );
  NOR21 U6988 ( .A(n6088), .B(n1828), .Q(n1811) );
  NOR21 U6989 ( .A(n6081), .B(n1790), .Q(n1776) );
  NOR21 U6990 ( .A(n1831), .B(n6090), .Q(n1853) );
  BUF2 U6991 ( .A(n6496), .Q(n6491) );
  INV3 U6992 ( .A(n5720), .Q(n6496) );
  BUF2 U6993 ( .A(n6502), .Q(n6497) );
  INV3 U6994 ( .A(n5719), .Q(n6502) );
  NOR21 U6995 ( .A(inst_out[24]), .B(n5723), .Q(n3370) );
  NOR21 U6996 ( .A(inst_out[19]), .B(n5724), .Q(n2702) );
  NOR21 U6997 ( .A(inst_out[16]), .B(n5726), .Q(n2688) );
  NOR21 U6998 ( .A(n5725), .B(n5727), .Q(n3355) );
  NOR21 U6999 ( .A(n5726), .B(n5728), .Q(n2687) );
  NOR21 U7000 ( .A(inst_out[21]), .B(n5727), .Q(n3356) );
  NOR21 U7001 ( .A(inst_out[18]), .B(n5728), .Q(n2690) );
  NOR21 U7002 ( .A(n5721), .B(n5723), .Q(n3354) );
  NOR21 U7003 ( .A(n5722), .B(n5724), .Q(n2686) );
  NOR21 U7004 ( .A(inst_out[17]), .B(n5722), .Q(n2689) );
  NOR21 U7005 ( .A(n1462), .B(n4287), .Q(n4286) );
  INV3 U7006 ( .A(n4289), .Q(n1462) );
  NAND22 U7007 ( .A(n3380), .B(n3381), .Q(n3377) );
  NAND22 U7008 ( .A(n3386), .B(n3387), .Q(n3383) );
  XNR21 U7009 ( .A(n1816), .B(pc_rom[15]), .Q(n1815) );
  XNR21 U7010 ( .A(n5716), .B(n5718), .Q(n1980) );
  NOR21 U7011 ( .A(n6086), .B(n5715), .Q(n1865) );
  NAND22 U7012 ( .A(n5715), .B(n6086), .Q(n1771) );
  XNR21 U7013 ( .A(n1781), .B(pc_rom[13]), .Q(n1779) );
  OAI311 U7014 ( .A(n1481), .B(n5699), .C(n5942), .D(n5700), .Q(n1854) );
  INV3 U7015 ( .A(rst), .Q(n1108) );
  CLKIN1 U7016 ( .A(n1768), .Q(n1255) );
  INV3 U7017 ( .A(n4333), .Q(n1414) );
  NOR21 U7018 ( .A(n4333), .B(n6761), .Q(n5812) );
  NAND31 U7019 ( .A(n1361), .B(n6199), .C(n1470), .Q(n3433) );
  NAND22 U7020 ( .A(n3436), .B(n6199), .Q(n3449) );
  INV3 U7021 ( .A(n6199), .Q(n1426) );
  INV0 U7022 ( .A(n4052), .Q(n1362) );
  NOR20 U7023 ( .A(n4227), .B(n6514), .Q(n4232) );
  NAND20 U7024 ( .A(n1470), .B(n4227), .Q(n4234) );
  INV3 U7025 ( .A(n4227), .Q(n1428) );
  OAI2112 U7026 ( .A(n6204), .B(n3692), .C(n3589), .D(n4247), .Q(n6264) );
  INV0 U7027 ( .A(n6280), .Q(n6266) );
  XNR21 U7028 ( .A(rs[4]), .B(n6268), .Q(n4555) );
  NAND30 U7029 ( .A(n5848), .B(n5941), .C(n5867), .Q(n6269) );
  NAND31 U7030 ( .A(\instruction_decode/old_ex [2]), .B(n1866), .C(
        \instruction_decode/old_ex [1]), .Q(n1841) );
  OAI211 U7031 ( .A(n6486), .B(n1157), .C(n1860), .Q(
        \instruction_fetch/pc_4 [7]) );
  OAI211 U7032 ( .A(n6487), .B(n5702), .C(n1829), .Q(n5794) );
  OAI211 U7033 ( .A(n5826), .B(n5703), .C(n1826), .Q(n5793) );
  OAI222 U7034 ( .A(n6308), .B(n6272), .C(n6288), .D(n6273), .Q(n6271) );
  XNR21 U7035 ( .A(pc_rom[28]), .B(n1853), .Q(n6273) );
  CLKIN3 U7036 ( .A(n6592), .Q(n6290) );
  CLKIN6 U7037 ( .A(n6311), .Q(n6287) );
  INV1 U7038 ( .A(n6313), .Q(n6274) );
  AOI220 U7039 ( .A(n1789), .B(n6311), .C(n1142), .D(inst_out[15]), .Q(n1788)
         );
  OAI220 U7040 ( .A(n6315), .B(n4579), .C(n6285), .D(n1850), .Q(n5801) );
  NOR20 U7041 ( .A(n6285), .B(n1138), .Q(n5764) );
  OAI220 U7042 ( .A(n6297), .B(n6276), .C(n6281), .D(n6277), .Q(n6275) );
  XNR21 U7043 ( .A(n4580), .B(n1864), .Q(n6277) );
  INV2 U7044 ( .A(n6592), .Q(n6289) );
  CLKIN3 U7045 ( .A(n6591), .Q(n6295) );
  CLKIN3 U7046 ( .A(n6591), .Q(n6296) );
  OAI211 U7047 ( .A(n5826), .B(n6262), .C(n1814), .Q(n5789) );
  OAI211 U7048 ( .A(n5826), .B(n5707), .C(n1788), .Q(n5778) );
  NOR21 U7049 ( .A(n6287), .B(n1120), .Q(n5746) );
  INV2 U7050 ( .A(n6307), .Q(n6300) );
  INV6 U7051 ( .A(n1780), .Q(n6310) );
  NOR20 U7052 ( .A(n1975), .B(n1976), .Q(\instruction_decode/old_ex [3]) );
  BUF2 U7053 ( .A(n1773), .Q(n6279) );
  OAI2110 U7054 ( .A(n5732), .B(n4406), .C(n5733), .D(n5699), .Q(n4405) );
  NAND20 U7055 ( .A(n5732), .B(n5733), .Q(n4412) );
  XNR20 U7056 ( .A(n5732), .B(n5999), .Q(n4416) );
  INV3 U7057 ( .A(n1967), .Q(n1146) );
  CLKIN1 U7058 ( .A(n6312), .Q(n6282) );
  CLKIN1 U7059 ( .A(n6283), .Q(n6285) );
  OAI221 U7060 ( .A(n4576), .B(n6298), .C(n6486), .D(n5709), .Q(n5781) );
  AOI220 U7061 ( .A(n6332), .B(data_2[23]), .C(n5815), .D(ram_adr[23]), .Q(
        n4442) );
  INV6 U7062 ( .A(n6311), .Q(n6286) );
  INV3 U7063 ( .A(n6289), .Q(n6291) );
  INV3 U7064 ( .A(n6290), .Q(n6294) );
  INV3 U7065 ( .A(n6591), .Q(n6297) );
  INV3 U7066 ( .A(n6297), .Q(n6302) );
  INV3 U7067 ( .A(n6297), .Q(n6303) );
  INV3 U7068 ( .A(n6287), .Q(n6304) );
  INV3 U7069 ( .A(n6304), .Q(n6305) );
  INV3 U7070 ( .A(n6304), .Q(n6306) );
  INV2 U7071 ( .A(n6278), .Q(n6315) );
  BUF2 U7072 ( .A(n6310), .Q(n6592) );
  BUF2 U7073 ( .A(n6310), .Q(n6591) );
  AOI221 U7074 ( .A(n1486), .B(ram_adr[3]), .C(n1484), .D(n6936), .Q(n4422) );
  NAND31 U7075 ( .A(n6513), .B(n4216), .C(n4172), .Q(n4230) );
  AOI210 U7076 ( .A(n4216), .B(n4217), .C(n4172), .Q(n4214) );
  NOR30 U7077 ( .A(n3407), .B(n4172), .C(n4216), .Q(n4226) );
  AOI210 U7078 ( .A(n4171), .B(n4170), .C(n4062), .Q(n4215) );
  XNR20 U7079 ( .A(rt[3]), .B(n5722), .Q(n3379) );
  XNR20 U7080 ( .A(rt[3]), .B(n5721), .Q(n3385) );
  XNR20 U7081 ( .A(write_register[3]), .B(rt[3]), .Q(n4560) );
  AOI2110 U7082 ( .A(n3949), .B(n3930), .C(n3950), .D(n1354), .Q(n3923) );
  OAI220 U7083 ( .A(n1284), .B(n3540), .C(n3930), .D(n3951), .Q(n3950) );
  OAI220 U7084 ( .A(n3930), .B(n3610), .C(n4333), .D(n3611), .Q(n4399) );
  OAI210 U7085 ( .A(n6204), .B(n3692), .C(n3690), .Q(n3935) );
  NOR40 U7086 ( .A(n5945), .B(n5868), .C(n6086), .D(n1974), .Q(
        \instruction_decode/old_ex [5]) );
  OAI220 U7087 ( .A(n3440), .B(n1362), .C(n4063), .D(n4062), .Q(n4140) );
  NOR31 U7088 ( .A(n3442), .B(n4062), .C(n4174), .Q(n4052) );
  OAI2110 U7089 ( .A(n1416), .B(n3685), .C(n3504), .D(n3686), .Q(n3679) );
  AOI310 U7090 ( .A(n3976), .B(n1308), .C(n6513), .D(n4043), .Q(n4042) );
  AOI310 U7091 ( .A(n6513), .B(n1308), .C(n4002), .D(n1348), .Q(n4040) );
  AOI220 U7092 ( .A(n6356), .B(n1416), .C(n1258), .D(n1414), .Q(n4371) );
  AOI220 U7093 ( .A(n6356), .B(n6347), .C(n1258), .D(n1416), .Q(n3702) );
  AOI210 U7094 ( .A(n1308), .B(n3913), .C(n3914), .Q(n3968) );
  OAI210 U7095 ( .A(n4024), .B(n1442), .C(n1308), .Q(n4000) );
  AOI220 U7096 ( .A(n1416), .B(n1294), .C(n6347), .D(n6353), .Q(n3945) );
  AOI220 U7097 ( .A(n4336), .B(n6349), .C(n1317), .D(n1416), .Q(n4330) );
  AOI220 U7098 ( .A(n1830), .B(n6315), .C(n1142), .D(n6497), .Q(n1829) );
  AOI220 U7099 ( .A(n6311), .B(n1815), .C(n1142), .D(inst_out[13]), .Q(n1814)
         );
  AOI220 U7100 ( .A(n1824), .B(n6313), .C(n1142), .D(inst_out[19]), .Q(n1823)
         );
  AOI220 U7101 ( .A(n1861), .B(n6312), .C(n1142), .D(inst_out[5]), .Q(n1860)
         );
  AOI220 U7102 ( .A(n1798), .B(n6312), .C(n1142), .D(inst_out[3]), .Q(n1797)
         );
  OAI210 U7103 ( .A(pc_out[2]), .B(n6311), .C(n6270), .Q(n1840) );
  AOI210 U7104 ( .A(n3589), .B(n3590), .C(n3591), .Q(n3588) );
  XNR20 U7105 ( .A(n6221), .B(n6317), .Q(n3376) );
  XNR20 U7106 ( .A(n6221), .B(n5719), .Q(n3382) );
  NAND30 U7107 ( .A(n3637), .B(n1386), .C(n3634), .Q(n3802) );
  XOR20 U7108 ( .A(rs[3]), .B(write_register_ex[3]), .Q(n4556) );
  OAI220 U7109 ( .A(n4577), .B(n6281), .C(n6486), .D(n5708), .Q(n5788) );
  OAI220 U7110 ( .A(n6267), .B(n5612), .C(n6992), .D(n6505), .Q(n4287) );
  NAND34 U7111 ( .A(n1308), .B(n3912), .C(n3913), .Q(n3634) );
  INV3 U7112 ( .A(n1867), .Q(n1147) );
  OAI210 U7113 ( .A(n5730), .B(n1973), .C(n1969), .Q(
        \instruction_decode/old_m [0]) );
  AOI2110 U7114 ( .A(n3537), .B(n3538), .C(n3539), .D(n1354), .Q(n3522) );
  OAI220 U7115 ( .A(n3538), .B(n6508), .C(n6348), .D(n6511), .Q(n3608) );
  OAI220 U7116 ( .A(n1283), .B(n3540), .C(n3538), .D(n3541), .Q(n3539) );
  OAI220 U7117 ( .A(n1420), .B(n6508), .C(n3538), .D(n6511), .Q(n3697) );
  AOI210 U7118 ( .A(n3561), .B(n1350), .C(n4050), .Q(n3440) );
  OAI220 U7119 ( .A(n3508), .B(n3477), .C(n3538), .D(n3542), .Q(n4327) );
  NAND31 U7120 ( .A(write_register[1]), .B(write_register[2]), .C(
        write_register[0]), .Q(n1961) );
  NAND31 U7121 ( .A(write_register[2]), .B(n5848), .C(write_register[0]), .Q(
        n1963) );
  NAND31 U7122 ( .A(write_register[1]), .B(n5941), .C(write_register[0]), .Q(
        n1957) );
  NAND31 U7123 ( .A(n5848), .B(n5941), .C(write_register[0]), .Q(n1959) );
  XNR20 U7124 ( .A(write_register[0]), .B(rs[0]), .Q(n4545) );
  XNR20 U7125 ( .A(n1485), .B(write_register[0]), .Q(n4564) );
  NAND28 U7126 ( .A(n1149), .B(n5730), .Q(n1975) );
  OAI220 U7127 ( .A(n1385), .B(n6352), .C(n6228), .D(n3617), .Q(n3987) );
  OAI220 U7128 ( .A(n1272), .B(n3540), .C(n6228), .D(n3682), .Q(n3680) );
  OAI220 U7129 ( .A(n6228), .B(n3610), .C(n3930), .D(n3611), .Q(n3929) );
  OAI220 U7130 ( .A(n6228), .B(n6508), .C(n1418), .D(n6511), .Q(n4398) );
  OAI220 U7131 ( .A(n1418), .B(n3610), .C(n6228), .D(n3611), .Q(n3698) );
  OAI210 U7132 ( .A(n3681), .B(n5817), .C(n3592), .Q(n4336) );
  AOI2110 U7133 ( .A(n1473), .B(n1461), .C(n6266), .D(n3620), .Q(n3619) );
  OAI220 U7134 ( .A(n1428), .B(n3404), .C(n4227), .D(n6517), .Q(n4225) );
  OAI310 U7135 ( .A(n3407), .B(n1296), .C(n4175), .D(n4234), .Q(n4233) );
  NOR21 U7136 ( .A(n4227), .B(n4176), .Q(n4320) );
  INV6 U7137 ( .A(n4041), .Q(n1308) );
  NAND30 U7138 ( .A(n6265), .B(data_2[3]), .C(n4424), .Q(n4421) );
  CLKBU15 U7139 ( .A(\execute/n459 ), .Q(n6349) );
endmodule

