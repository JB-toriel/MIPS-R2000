//-----------------------------------------------------
	// This is design of the fetch stage of the pipeline
	// Design Name : IF
	// File Name   : fetch.sv
	// Function    :
	// Authors     : de Sainte Marie Nils - Edde Jean-Baptiste
//-----------------------------------------------------

/*
module NOM (LISTE DES PORTS);

DECLARATION DES PORTS
DECLARATION DES PARAMETRES

`include "NOM DE FICHIER";

DECLARATIONS DE VARIABLES
AFFECTATIONS
INSTANCIATIONS DE SOUS-MODULES
BLOCS initial ET always
TACHES ET FONCTIONS

endmodule
*/

/*
	Inputs : internally must always be of type net, externally the inputs can be connected to a variable of type reg or net.
	Outputs : internally can be of type net or reg, externally the outputs must be connected to a variable of type net.
	Inouts : internally or externally must always be type net, can only be connected to a variable net type.
*/


module ID ( inst_in, inst_2521, inst_2016, inst_1511/*, ...*/);
	input [31:0] inst_in;
	output reg [4:0] inst_2521, inst_2016, inst_1511;

  	always@(inst_in)
  		begin
          inst_2521 <= inst_in[25:21];
          inst_2016 <= inst_in[20:16];
          inst_1511 <= inst_in[15:11];
        end

	endmodule // End of ID module
